`define HLS_NAME DigitRec
