`define HLS_NAME face_detect
