module axis_fifo_wrapper_losscheck #
(
  parameter ASSERT_ON = 1'b1
)
(
  input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [31:0] s_axis_tdata,
  input logic [3:0] s_axis_tkeep,
  input logic [0:0] s_axis_tvalid,
  output logic [0:0] s_axis_tready,
  input logic [0:0] s_axis_tlast,
  input logic [0:0] s_axis_tuser,
  output logic [31:0] m_axis_tdata,
  output logic [3:0] m_axis_tkeep,
  output logic [0:0] m_axis_tvalid,
  input logic [0:0] m_axis_tready,
  output logic [0:0] m_axis_tlast,
  output logic [0:0] m_axis_tuser,
  output logic [0:0] status_overflow,
  output logic [0:0] status_bad_frame,
  output logic [0:0] status_good_frame,
  output logic [0:0] status_empty
);

  logic [63:0] TASKPASS_cycle_counter ;
  logic [10:0] axis_fifo_inst__DOT__wr_ptr_reg ;
  logic [10:0] axis_fifo_inst__DOT__wr_ptr_next ;
  logic [10:0] axis_fifo_inst__DOT__wr_ptr_cur_reg ;
  logic [10:0] axis_fifo_inst__DOT__wr_ptr_cur_next ;
  logic [10:0] axis_fifo_inst__DOT__wr_addr_reg ;
  logic [10:0] axis_fifo_inst__DOT__rd_ptr_reg ;
  logic [10:0] axis_fifo_inst__DOT__rd_ptr_next ;
  logic [10:0] axis_fifo_inst__DOT__rd_addr_reg ;
  logic [37:0] axis_fifo_inst__DOT__mem [1023:0] ;
  logic [37:0] axis_fifo_inst__DOT__mem_read_data_reg ;
  logic [0:0] axis_fifo_inst__DOT__mem_read_data_valid_reg ;
  logic [0:0] axis_fifo_inst__DOT__mem_read_data_valid_next ;
  logic [37:0] axis_fifo_inst__DOT__s_axis ;
  logic [37:0] axis_fifo_inst__DOT__m_axis_reg ;
  logic [0:0] axis_fifo_inst__DOT__m_axis_tvalid_reg ;
  logic [0:0] axis_fifo_inst__DOT__m_axis_tvalid_next ;
  logic [0:0] axis_fifo_inst__DOT__full ;
  logic [0:0] axis_fifo_inst__DOT__empty ;
  logic [0:0] axis_fifo_inst__DOT__full_cur ;
  logic [0:0] axis_fifo_inst__DOT__write ;
  logic [0:0] axis_fifo_inst__DOT__read ;
  logic [0:0] axis_fifo_inst__DOT__store_output ;
  logic [0:0] axis_fifo_inst__DOT__drop_frame_reg ;
  logic [0:0] axis_fifo_inst__DOT__drop_frame_next ;
  logic [0:0] axis_fifo_inst__DOT__overflow_reg ;
  logic [0:0] axis_fifo_inst__DOT__overflow_next ;
  logic [0:0] axis_fifo_inst__DOT__bad_frame_reg ;
  logic [0:0] axis_fifo_inst__DOT__bad_frame_next ;
  logic [0:0] axis_fifo_inst__DOT__good_frame_reg ;
  logic [0:0] axis_fifo_inst__DOT__good_frame_next ;
  assign axis_fifo_inst__DOT__full = (axis_fifo_inst__DOT__wr_ptr_reg[10] != axis_fifo_inst__DOT__rd_ptr_reg[10]) & (axis_fifo_inst__DOT__wr_ptr_reg[9:0] == axis_fifo_inst__DOT__rd_ptr_reg[9:0]);
  assign axis_fifo_inst__DOT__empty = axis_fifo_inst__DOT__wr_ptr_reg == axis_fifo_inst__DOT__rd_ptr_reg;
  assign status_empty = axis_fifo_inst__DOT__empty;
  assign axis_fifo_inst__DOT__full_cur = (axis_fifo_inst__DOT__wr_ptr_reg[10] != axis_fifo_inst__DOT__wr_ptr_cur_reg[10]) & (axis_fifo_inst__DOT__wr_ptr_reg[9:0] == axis_fifo_inst__DOT__wr_ptr_cur_reg[9:0]);
  assign s_axis_tready = ~axis_fifo_inst__DOT__full;
  assign axis_fifo_inst__DOT__s_axis[31:0] = s_axis_tdata;
  assign axis_fifo_inst__DOT__s_axis[35:32] = s_axis_tkeep;
  assign axis_fifo_inst__DOT__s_axis[36] = s_axis_tlast;
  assign axis_fifo_inst__DOT__s_axis[37] = s_axis_tuser;
  assign m_axis_tvalid = axis_fifo_inst__DOT__m_axis_tvalid_reg;
  assign m_axis_tdata = axis_fifo_inst__DOT__m_axis_reg[31:0];
  assign m_axis_tkeep = axis_fifo_inst__DOT__m_axis_reg[35:32];
  assign m_axis_tlast = axis_fifo_inst__DOT__m_axis_reg[36];
  assign m_axis_tuser = axis_fifo_inst__DOT__m_axis_reg[37];
  assign status_overflow = axis_fifo_inst__DOT__overflow_reg;
  assign status_bad_frame = axis_fifo_inst__DOT__bad_frame_reg;
  assign status_good_frame = axis_fifo_inst__DOT__good_frame_reg;

  always_comb begin
    axis_fifo_inst__DOT__write = 1'h0;
    axis_fifo_inst__DOT__drop_frame_next = 1'h0;
    axis_fifo_inst__DOT__overflow_next = 1'h0;
    axis_fifo_inst__DOT__bad_frame_next = 1'h0;
    axis_fifo_inst__DOT__good_frame_next = 1'h0;
    axis_fifo_inst__DOT__wr_ptr_next = axis_fifo_inst__DOT__wr_ptr_reg;
    axis_fifo_inst__DOT__wr_ptr_cur_next = axis_fifo_inst__DOT__wr_ptr_cur_reg;
    if (s_axis_tvalid) begin
      if (~axis_fifo_inst__DOT__full) begin
        if (axis_fifo_inst__DOT__full | axis_fifo_inst__DOT__full_cur | axis_fifo_inst__DOT__drop_frame_reg) begin
          axis_fifo_inst__DOT__drop_frame_next = 1'h1;
          if (s_axis_tlast) begin
            axis_fifo_inst__DOT__wr_ptr_cur_next = axis_fifo_inst__DOT__wr_ptr_reg;
            axis_fifo_inst__DOT__drop_frame_next = 1'h0;
            axis_fifo_inst__DOT__overflow_next = 1'h1;
          end 
        end else begin
          axis_fifo_inst__DOT__write = 1'h1;
          axis_fifo_inst__DOT__wr_ptr_cur_next = 11'h1 + axis_fifo_inst__DOT__wr_ptr_cur_reg;
          if (s_axis_tlast) begin
            axis_fifo_inst__DOT__wr_ptr_next = 11'h1 + axis_fifo_inst__DOT__wr_ptr_cur_reg;
            axis_fifo_inst__DOT__good_frame_next = 1'h1;
          end 
        end
      end 
    end 
  end

  always_comb begin
    axis_fifo_inst__DOT__read = 1'h0;
    axis_fifo_inst__DOT__rd_ptr_next = axis_fifo_inst__DOT__rd_ptr_reg;
    axis_fifo_inst__DOT__mem_read_data_valid_next = axis_fifo_inst__DOT__mem_read_data_valid_reg;
    if (axis_fifo_inst__DOT__store_output | ~axis_fifo_inst__DOT__mem_read_data_valid_reg) begin
      if (axis_fifo_inst__DOT__empty) begin
        axis_fifo_inst__DOT__mem_read_data_valid_next = 1'h0;
      end else begin
        axis_fifo_inst__DOT__read = 1'h1;
        axis_fifo_inst__DOT__mem_read_data_valid_next = 1'h1;
        axis_fifo_inst__DOT__rd_ptr_next = 11'h1 + axis_fifo_inst__DOT__rd_ptr_reg;
      end
    end 
  end

  always_comb begin
    axis_fifo_inst__DOT__store_output = 1'h0;
    axis_fifo_inst__DOT__m_axis_tvalid_next = axis_fifo_inst__DOT__m_axis_tvalid_reg;
    if (m_axis_tready | ~m_axis_tvalid) begin
      axis_fifo_inst__DOT__store_output = 1'h1;
      axis_fifo_inst__DOT__m_axis_tvalid_next = axis_fifo_inst__DOT__mem_read_data_valid_reg;
    end 
  end

  initial begin
    axis_fifo_inst__DOT__wr_ptr_reg = 11'h0;
    axis_fifo_inst__DOT__wr_ptr_cur_reg = 11'h0;
    axis_fifo_inst__DOT__wr_addr_reg = 11'h0;
    axis_fifo_inst__DOT__rd_ptr_reg = 11'h0;
    axis_fifo_inst__DOT__rd_addr_reg = 11'h0;
    axis_fifo_inst__DOT__mem_read_data_valid_reg = 1'h0;
    axis_fifo_inst__DOT__m_axis_tvalid_reg = 1'h0;
    axis_fifo_inst__DOT__drop_frame_reg = 1'h0;
    axis_fifo_inst__DOT__overflow_reg = 1'h0;
    axis_fifo_inst__DOT__bad_frame_reg = 1'h0;
    axis_fifo_inst__DOT__good_frame_reg = 1'h0;
  end

  always @(posedge clk) begin
    if (rst) begin
      axis_fifo_inst__DOT__wr_ptr_reg <= 11'h0;
      axis_fifo_inst__DOT__wr_ptr_cur_reg <= 11'h0;
      axis_fifo_inst__DOT__drop_frame_reg <= 1'h0;
      axis_fifo_inst__DOT__overflow_reg <= 1'h0;
      axis_fifo_inst__DOT__bad_frame_reg <= 1'h0;
      axis_fifo_inst__DOT__good_frame_reg <= 1'h0;
    end else begin
      axis_fifo_inst__DOT__wr_ptr_reg <= axis_fifo_inst__DOT__wr_ptr_next;
      axis_fifo_inst__DOT__wr_ptr_cur_reg <= axis_fifo_inst__DOT__wr_ptr_cur_next;
      axis_fifo_inst__DOT__drop_frame_reg <= axis_fifo_inst__DOT__drop_frame_next;
      axis_fifo_inst__DOT__overflow_reg <= axis_fifo_inst__DOT__overflow_next;
      axis_fifo_inst__DOT__bad_frame_reg <= axis_fifo_inst__DOT__bad_frame_next;
      axis_fifo_inst__DOT__good_frame_reg <= axis_fifo_inst__DOT__good_frame_next;
    end
    axis_fifo_inst__DOT__wr_addr_reg <= axis_fifo_inst__DOT__wr_ptr_cur_next;
    if (axis_fifo_inst__DOT__write) begin
      axis_fifo_inst__DOT__mem[axis_fifo_inst__DOT__wr_addr_reg[9:0]] <= axis_fifo_inst__DOT__s_axis;
    end 
  end

  always @(posedge clk) begin
    if (rst) begin
      axis_fifo_inst__DOT__rd_ptr_reg <= 11'h0;
      axis_fifo_inst__DOT__mem_read_data_valid_reg <= 1'h0;
    end else begin
      axis_fifo_inst__DOT__rd_ptr_reg <= axis_fifo_inst__DOT__rd_ptr_next;
      axis_fifo_inst__DOT__mem_read_data_valid_reg <= axis_fifo_inst__DOT__mem_read_data_valid_next;
    end
    axis_fifo_inst__DOT__rd_addr_reg <= axis_fifo_inst__DOT__rd_ptr_next;
    if (axis_fifo_inst__DOT__read) begin
      axis_fifo_inst__DOT__mem_read_data_reg <= axis_fifo_inst__DOT__mem[axis_fifo_inst__DOT__rd_addr_reg[9:0]];
    end 
  end

  always @(posedge clk) begin
    axis_fifo_inst__DOT__m_axis_tvalid_reg <= ~rst & axis_fifo_inst__DOT__m_axis_tvalid_next;
    if (axis_fifo_inst__DOT__store_output) begin
      axis_fifo_inst__DOT__m_axis_reg <= axis_fifo_inst__DOT__mem_read_data_reg;
    end 
  end
  logic m_axis_tdata__BRA__31__03A0__KET____AV__ ;
  logic m_axis_tdata__BRA__31__03A0__KET____AI__ ;
  logic m_axis_tdata__BRA__31__03A0__KET____ASSIGN__ ;
  logic m_axis_tdata__BRA__31__03A0__KET____VALID__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AI__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____ASSIGN__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____VALID__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV_Q__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AI_Q__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____ASSIGN_Q__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____VALID_Q__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AI__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____VALID__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV_Q__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AI_Q__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN_Q__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____VALID_Q__ ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__ [1023:0] ;
  logic axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____AV__ ;
  logic axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____AI__ ;
  logic axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____ASSIGN__ ;
  logic axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____PROP__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____PROP_Q__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____GOOD__ ;
  logic axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____GOOD_Q__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP_Q__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD__ ;
  logic axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD_Q__ ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__ [1023:0] ;
  logic axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__ [1023:0] ;
  logic [9:0] array_pointer_delay_0 ;
  logic s_axis_tdata__VALID__ ;
  assign m_axis_tdata__BRA__31__03A0__KET____AV__ = axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____VALID__;
  assign m_axis_tdata__BRA__31__03A0__KET____AI__ = m_axis_tdata__BRA__31__03A0__KET____ASSIGN__ & ~m_axis_tdata__BRA__31__03A0__KET____AV__;
  assign m_axis_tdata__BRA__31__03A0__KET____ASSIGN__ = 1'b1;
  assign m_axis_tdata__BRA__31__03A0__KET____VALID__ = m_axis_tdata__BRA__31__03A0__KET____AV__;
  assign axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV__ = axis_fifo_inst__DOT__store_output & axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____VALID__;
  assign axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AI__ = axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____ASSIGN__ & ~axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV__;
  assign axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____ASSIGN__ = axis_fifo_inst__DOT__store_output;
  assign axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____VALID__ = axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV_Q__ | ~axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____ASSIGN_Q__ & axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____VALID_Q__;
  assign axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV__ = axis_fifo_inst__DOT__read & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[axis_fifo_inst__DOT__rd_addr_reg[9:0]];
  assign axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AI__ = axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN__ & ~axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV__;
  assign axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN__ = axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____VALID__ = axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV_Q__ | ~axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN_Q__ & axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____VALID_Q__;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h0] = (10'h0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h0] = axis_fifo_inst__DOT__write & (10'h0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1] = (10'h1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1] = axis_fifo_inst__DOT__write & (10'h1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2] = (10'h2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2] = axis_fifo_inst__DOT__write & (10'h2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3] = (10'h3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3] = axis_fifo_inst__DOT__write & (10'h3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4] = (10'h4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4] = axis_fifo_inst__DOT__write & (10'h4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5] = (10'h5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5] = axis_fifo_inst__DOT__write & (10'h5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6] = (10'h6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6] = axis_fifo_inst__DOT__write & (10'h6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7] = (10'h7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7] = axis_fifo_inst__DOT__write & (10'h7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8] = (10'h8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8] = axis_fifo_inst__DOT__write & (10'h8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9] = (10'h9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9] = axis_fifo_inst__DOT__write & (10'h9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha] = (10'ha == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha] = axis_fifo_inst__DOT__write & (10'ha == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb] = (10'hb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb] = axis_fifo_inst__DOT__write & (10'hb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc] = (10'hc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc] = axis_fifo_inst__DOT__write & (10'hc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd] = (10'hd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd] = axis_fifo_inst__DOT__write & (10'hd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he] = (10'he == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he] = axis_fifo_inst__DOT__write & (10'he == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf] = (10'hf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf] = axis_fifo_inst__DOT__write & (10'hf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10] = (10'h10 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10] = axis_fifo_inst__DOT__write & (10'h10 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11] = (10'h11 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11] = axis_fifo_inst__DOT__write & (10'h11 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12] = (10'h12 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12] = axis_fifo_inst__DOT__write & (10'h12 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13] = (10'h13 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13] = axis_fifo_inst__DOT__write & (10'h13 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14] = (10'h14 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14] = axis_fifo_inst__DOT__write & (10'h14 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15] = (10'h15 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15] = axis_fifo_inst__DOT__write & (10'h15 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16] = (10'h16 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16] = axis_fifo_inst__DOT__write & (10'h16 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17] = (10'h17 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17] = axis_fifo_inst__DOT__write & (10'h17 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18] = (10'h18 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18] = axis_fifo_inst__DOT__write & (10'h18 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19] = (10'h19 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19] = axis_fifo_inst__DOT__write & (10'h19 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a] = (10'h1a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a] = axis_fifo_inst__DOT__write & (10'h1a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b] = (10'h1b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b] = axis_fifo_inst__DOT__write & (10'h1b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c] = (10'h1c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c] = axis_fifo_inst__DOT__write & (10'h1c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d] = (10'h1d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d] = axis_fifo_inst__DOT__write & (10'h1d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e] = (10'h1e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e] = axis_fifo_inst__DOT__write & (10'h1e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f] = (10'h1f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f] = axis_fifo_inst__DOT__write & (10'h1f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20] = (10'h20 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20] = axis_fifo_inst__DOT__write & (10'h20 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21] = (10'h21 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21] = axis_fifo_inst__DOT__write & (10'h21 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22] = (10'h22 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22] = axis_fifo_inst__DOT__write & (10'h22 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23] = (10'h23 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23] = axis_fifo_inst__DOT__write & (10'h23 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24] = (10'h24 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24] = axis_fifo_inst__DOT__write & (10'h24 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25] = (10'h25 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25] = axis_fifo_inst__DOT__write & (10'h25 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26] = (10'h26 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26] = axis_fifo_inst__DOT__write & (10'h26 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27] = (10'h27 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27] = axis_fifo_inst__DOT__write & (10'h27 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28] = (10'h28 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28] = axis_fifo_inst__DOT__write & (10'h28 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29] = (10'h29 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29] = axis_fifo_inst__DOT__write & (10'h29 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a] = (10'h2a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a] = axis_fifo_inst__DOT__write & (10'h2a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b] = (10'h2b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b] = axis_fifo_inst__DOT__write & (10'h2b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c] = (10'h2c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c] = axis_fifo_inst__DOT__write & (10'h2c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d] = (10'h2d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d] = axis_fifo_inst__DOT__write & (10'h2d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e] = (10'h2e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e] = axis_fifo_inst__DOT__write & (10'h2e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f] = (10'h2f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f] = axis_fifo_inst__DOT__write & (10'h2f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30] = (10'h30 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30] = axis_fifo_inst__DOT__write & (10'h30 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31] = (10'h31 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31] = axis_fifo_inst__DOT__write & (10'h31 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32] = (10'h32 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32] = axis_fifo_inst__DOT__write & (10'h32 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33] = (10'h33 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33] = axis_fifo_inst__DOT__write & (10'h33 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34] = (10'h34 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34] = axis_fifo_inst__DOT__write & (10'h34 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35] = (10'h35 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35] = axis_fifo_inst__DOT__write & (10'h35 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36] = (10'h36 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36] = axis_fifo_inst__DOT__write & (10'h36 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37] = (10'h37 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37] = axis_fifo_inst__DOT__write & (10'h37 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38] = (10'h38 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38] = axis_fifo_inst__DOT__write & (10'h38 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39] = (10'h39 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39] = axis_fifo_inst__DOT__write & (10'h39 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a] = (10'h3a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a] = axis_fifo_inst__DOT__write & (10'h3a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b] = (10'h3b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b] = axis_fifo_inst__DOT__write & (10'h3b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c] = (10'h3c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c] = axis_fifo_inst__DOT__write & (10'h3c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d] = (10'h3d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d] = axis_fifo_inst__DOT__write & (10'h3d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e] = (10'h3e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e] = axis_fifo_inst__DOT__write & (10'h3e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f] = (10'h3f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f] = axis_fifo_inst__DOT__write & (10'h3f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h40] = (10'h40 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h40] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h40] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h40];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h40] = axis_fifo_inst__DOT__write & (10'h40 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h40] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h40] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h40] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h40];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h41] = (10'h41 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h41] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h41] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h41];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h41] = axis_fifo_inst__DOT__write & (10'h41 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h41] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h41] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h41] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h41];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h42] = (10'h42 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h42] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h42] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h42];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h42] = axis_fifo_inst__DOT__write & (10'h42 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h42] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h42] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h42] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h42];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h43] = (10'h43 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h43] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h43] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h43];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h43] = axis_fifo_inst__DOT__write & (10'h43 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h43] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h43] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h43] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h43];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h44] = (10'h44 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h44] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h44] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h44];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h44] = axis_fifo_inst__DOT__write & (10'h44 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h44] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h44] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h44] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h44];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h45] = (10'h45 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h45] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h45] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h45];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h45] = axis_fifo_inst__DOT__write & (10'h45 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h45] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h45] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h45] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h45];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h46] = (10'h46 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h46] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h46] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h46];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h46] = axis_fifo_inst__DOT__write & (10'h46 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h46] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h46] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h46] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h46];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h47] = (10'h47 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h47] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h47] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h47];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h47] = axis_fifo_inst__DOT__write & (10'h47 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h47] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h47] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h47] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h47];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h48] = (10'h48 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h48] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h48] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h48];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h48] = axis_fifo_inst__DOT__write & (10'h48 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h48] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h48] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h48] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h48];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h49] = (10'h49 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h49] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h49] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h49];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h49] = axis_fifo_inst__DOT__write & (10'h49 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h49] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h49] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h49] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h49];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4a] = (10'h4a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4a] = axis_fifo_inst__DOT__write & (10'h4a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4b] = (10'h4b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4b] = axis_fifo_inst__DOT__write & (10'h4b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4c] = (10'h4c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4c] = axis_fifo_inst__DOT__write & (10'h4c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4d] = (10'h4d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4d] = axis_fifo_inst__DOT__write & (10'h4d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4e] = (10'h4e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4e] = axis_fifo_inst__DOT__write & (10'h4e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4f] = (10'h4f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4f] = axis_fifo_inst__DOT__write & (10'h4f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h50] = (10'h50 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h50] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h50] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h50];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h50] = axis_fifo_inst__DOT__write & (10'h50 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h50] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h50] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h50] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h50];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h51] = (10'h51 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h51] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h51] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h51];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h51] = axis_fifo_inst__DOT__write & (10'h51 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h51] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h51] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h51] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h51];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h52] = (10'h52 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h52] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h52] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h52];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h52] = axis_fifo_inst__DOT__write & (10'h52 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h52] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h52] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h52] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h52];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h53] = (10'h53 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h53] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h53] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h53];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h53] = axis_fifo_inst__DOT__write & (10'h53 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h53] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h53] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h53] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h53];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h54] = (10'h54 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h54] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h54] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h54];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h54] = axis_fifo_inst__DOT__write & (10'h54 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h54] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h54] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h54] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h54];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h55] = (10'h55 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h55] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h55] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h55];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h55] = axis_fifo_inst__DOT__write & (10'h55 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h55] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h55] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h55] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h55];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h56] = (10'h56 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h56] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h56] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h56];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h56] = axis_fifo_inst__DOT__write & (10'h56 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h56] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h56] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h56] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h56];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h57] = (10'h57 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h57] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h57] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h57];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h57] = axis_fifo_inst__DOT__write & (10'h57 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h57] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h57] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h57] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h57];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h58] = (10'h58 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h58] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h58] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h58];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h58] = axis_fifo_inst__DOT__write & (10'h58 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h58] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h58] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h58] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h58];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h59] = (10'h59 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h59] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h59] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h59];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h59] = axis_fifo_inst__DOT__write & (10'h59 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h59] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h59] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h59] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h59];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5a] = (10'h5a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5a] = axis_fifo_inst__DOT__write & (10'h5a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5b] = (10'h5b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5b] = axis_fifo_inst__DOT__write & (10'h5b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5c] = (10'h5c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5c] = axis_fifo_inst__DOT__write & (10'h5c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5d] = (10'h5d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5d] = axis_fifo_inst__DOT__write & (10'h5d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5e] = (10'h5e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5e] = axis_fifo_inst__DOT__write & (10'h5e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5f] = (10'h5f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5f] = axis_fifo_inst__DOT__write & (10'h5f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h60] = (10'h60 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h60] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h60] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h60];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h60] = axis_fifo_inst__DOT__write & (10'h60 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h60] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h60] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h60] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h60];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h61] = (10'h61 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h61] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h61] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h61];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h61] = axis_fifo_inst__DOT__write & (10'h61 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h61] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h61] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h61] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h61];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h62] = (10'h62 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h62] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h62] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h62];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h62] = axis_fifo_inst__DOT__write & (10'h62 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h62] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h62] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h62] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h62];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h63] = (10'h63 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h63] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h63] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h63];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h63] = axis_fifo_inst__DOT__write & (10'h63 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h63] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h63] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h63] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h63];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h64] = (10'h64 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h64] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h64] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h64];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h64] = axis_fifo_inst__DOT__write & (10'h64 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h64] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h64] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h64] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h64];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h65] = (10'h65 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h65] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h65] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h65];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h65] = axis_fifo_inst__DOT__write & (10'h65 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h65] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h65] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h65] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h65];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h66] = (10'h66 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h66] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h66] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h66];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h66] = axis_fifo_inst__DOT__write & (10'h66 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h66] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h66] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h66] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h66];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h67] = (10'h67 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h67] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h67] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h67];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h67] = axis_fifo_inst__DOT__write & (10'h67 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h67] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h67] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h67] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h67];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h68] = (10'h68 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h68] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h68] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h68];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h68] = axis_fifo_inst__DOT__write & (10'h68 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h68] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h68] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h68] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h68];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h69] = (10'h69 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h69] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h69] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h69];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h69] = axis_fifo_inst__DOT__write & (10'h69 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h69] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h69] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h69] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h69];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6a] = (10'h6a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6a] = axis_fifo_inst__DOT__write & (10'h6a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6b] = (10'h6b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6b] = axis_fifo_inst__DOT__write & (10'h6b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6c] = (10'h6c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6c] = axis_fifo_inst__DOT__write & (10'h6c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6d] = (10'h6d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6d] = axis_fifo_inst__DOT__write & (10'h6d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6e] = (10'h6e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6e] = axis_fifo_inst__DOT__write & (10'h6e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6f] = (10'h6f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6f] = axis_fifo_inst__DOT__write & (10'h6f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h70] = (10'h70 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h70] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h70] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h70];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h70] = axis_fifo_inst__DOT__write & (10'h70 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h70] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h70] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h70] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h70];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h71] = (10'h71 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h71] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h71] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h71];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h71] = axis_fifo_inst__DOT__write & (10'h71 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h71] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h71] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h71] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h71];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h72] = (10'h72 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h72] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h72] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h72];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h72] = axis_fifo_inst__DOT__write & (10'h72 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h72] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h72] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h72] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h72];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h73] = (10'h73 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h73] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h73] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h73];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h73] = axis_fifo_inst__DOT__write & (10'h73 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h73] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h73] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h73] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h73];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h74] = (10'h74 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h74] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h74] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h74];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h74] = axis_fifo_inst__DOT__write & (10'h74 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h74] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h74] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h74] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h74];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h75] = (10'h75 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h75] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h75] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h75];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h75] = axis_fifo_inst__DOT__write & (10'h75 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h75] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h75] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h75] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h75];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h76] = (10'h76 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h76] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h76] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h76];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h76] = axis_fifo_inst__DOT__write & (10'h76 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h76] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h76] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h76] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h76];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h77] = (10'h77 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h77] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h77] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h77];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h77] = axis_fifo_inst__DOT__write & (10'h77 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h77] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h77] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h77] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h77];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h78] = (10'h78 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h78] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h78] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h78];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h78] = axis_fifo_inst__DOT__write & (10'h78 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h78] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h78] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h78] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h78];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h79] = (10'h79 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h79] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h79] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h79];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h79] = axis_fifo_inst__DOT__write & (10'h79 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h79] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h79] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h79] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h79];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7a] = (10'h7a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7a] = axis_fifo_inst__DOT__write & (10'h7a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7b] = (10'h7b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7b] = axis_fifo_inst__DOT__write & (10'h7b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7c] = (10'h7c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7c] = axis_fifo_inst__DOT__write & (10'h7c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7d] = (10'h7d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7d] = axis_fifo_inst__DOT__write & (10'h7d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7e] = (10'h7e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7e] = axis_fifo_inst__DOT__write & (10'h7e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7f] = (10'h7f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7f] = axis_fifo_inst__DOT__write & (10'h7f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h80] = (10'h80 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h80] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h80] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h80];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h80] = axis_fifo_inst__DOT__write & (10'h80 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h80] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h80] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h80] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h80];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h81] = (10'h81 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h81] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h81] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h81];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h81] = axis_fifo_inst__DOT__write & (10'h81 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h81] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h81] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h81] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h81];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h82] = (10'h82 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h82] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h82] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h82];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h82] = axis_fifo_inst__DOT__write & (10'h82 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h82] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h82] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h82] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h82];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h83] = (10'h83 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h83] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h83] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h83];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h83] = axis_fifo_inst__DOT__write & (10'h83 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h83] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h83] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h83] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h83];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h84] = (10'h84 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h84] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h84] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h84];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h84] = axis_fifo_inst__DOT__write & (10'h84 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h84] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h84] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h84] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h84];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h85] = (10'h85 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h85] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h85] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h85];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h85] = axis_fifo_inst__DOT__write & (10'h85 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h85] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h85] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h85] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h85];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h86] = (10'h86 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h86] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h86] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h86];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h86] = axis_fifo_inst__DOT__write & (10'h86 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h86] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h86] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h86] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h86];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h87] = (10'h87 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h87] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h87] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h87];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h87] = axis_fifo_inst__DOT__write & (10'h87 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h87] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h87] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h87] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h87];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h88] = (10'h88 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h88] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h88] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h88];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h88] = axis_fifo_inst__DOT__write & (10'h88 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h88] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h88] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h88] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h88];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h89] = (10'h89 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h89] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h89] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h89];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h89] = axis_fifo_inst__DOT__write & (10'h89 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h89] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h89] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h89] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h89];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8a] = (10'h8a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8a] = axis_fifo_inst__DOT__write & (10'h8a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8b] = (10'h8b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8b] = axis_fifo_inst__DOT__write & (10'h8b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8c] = (10'h8c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8c] = axis_fifo_inst__DOT__write & (10'h8c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8d] = (10'h8d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8d] = axis_fifo_inst__DOT__write & (10'h8d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8e] = (10'h8e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8e] = axis_fifo_inst__DOT__write & (10'h8e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8f] = (10'h8f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8f] = axis_fifo_inst__DOT__write & (10'h8f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h90] = (10'h90 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h90] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h90] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h90];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h90] = axis_fifo_inst__DOT__write & (10'h90 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h90] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h90] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h90] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h90];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h91] = (10'h91 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h91] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h91] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h91];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h91] = axis_fifo_inst__DOT__write & (10'h91 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h91] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h91] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h91] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h91];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h92] = (10'h92 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h92] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h92] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h92];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h92] = axis_fifo_inst__DOT__write & (10'h92 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h92] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h92] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h92] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h92];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h93] = (10'h93 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h93] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h93] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h93];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h93] = axis_fifo_inst__DOT__write & (10'h93 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h93] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h93] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h93] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h93];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h94] = (10'h94 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h94] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h94] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h94];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h94] = axis_fifo_inst__DOT__write & (10'h94 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h94] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h94] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h94] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h94];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h95] = (10'h95 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h95] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h95] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h95];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h95] = axis_fifo_inst__DOT__write & (10'h95 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h95] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h95] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h95] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h95];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h96] = (10'h96 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h96] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h96] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h96];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h96] = axis_fifo_inst__DOT__write & (10'h96 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h96] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h96] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h96] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h96];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h97] = (10'h97 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h97] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h97] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h97];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h97] = axis_fifo_inst__DOT__write & (10'h97 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h97] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h97] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h97] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h97];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h98] = (10'h98 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h98] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h98] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h98];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h98] = axis_fifo_inst__DOT__write & (10'h98 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h98] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h98] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h98] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h98];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h99] = (10'h99 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h99] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h99] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h99];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h99] = axis_fifo_inst__DOT__write & (10'h99 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h99] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h99] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h99] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h99];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9a] = (10'h9a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9a] = axis_fifo_inst__DOT__write & (10'h9a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9b] = (10'h9b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9b] = axis_fifo_inst__DOT__write & (10'h9b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9c] = (10'h9c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9c] = axis_fifo_inst__DOT__write & (10'h9c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9d] = (10'h9d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9d] = axis_fifo_inst__DOT__write & (10'h9d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9e] = (10'h9e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9e] = axis_fifo_inst__DOT__write & (10'h9e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9f] = (10'h9f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9f] = axis_fifo_inst__DOT__write & (10'h9f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha0] = (10'ha0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha0] = axis_fifo_inst__DOT__write & (10'ha0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha1] = (10'ha1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha1] = axis_fifo_inst__DOT__write & (10'ha1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha2] = (10'ha2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha2] = axis_fifo_inst__DOT__write & (10'ha2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha3] = (10'ha3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha3] = axis_fifo_inst__DOT__write & (10'ha3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha4] = (10'ha4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha4] = axis_fifo_inst__DOT__write & (10'ha4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha5] = (10'ha5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha5] = axis_fifo_inst__DOT__write & (10'ha5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha6] = (10'ha6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha6] = axis_fifo_inst__DOT__write & (10'ha6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha7] = (10'ha7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha7] = axis_fifo_inst__DOT__write & (10'ha7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha8] = (10'ha8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha8] = axis_fifo_inst__DOT__write & (10'ha8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha9] = (10'ha9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha9] = axis_fifo_inst__DOT__write & (10'ha9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'haa] = (10'haa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'haa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'haa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'haa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'haa] = axis_fifo_inst__DOT__write & (10'haa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'haa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'haa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'haa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'haa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hab] = (10'hab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hab] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hab] = axis_fifo_inst__DOT__write & (10'hab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hab] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hab] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hac] = (10'hac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hac] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hac] = axis_fifo_inst__DOT__write & (10'hac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hac] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hac] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'had] = (10'had == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'had] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'had] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'had];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'had] = axis_fifo_inst__DOT__write & (10'had == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'had] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'had] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'had] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'had];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hae] = (10'hae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hae] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hae] = axis_fifo_inst__DOT__write & (10'hae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hae] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hae] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'haf] = (10'haf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'haf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'haf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'haf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'haf] = axis_fifo_inst__DOT__write & (10'haf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'haf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'haf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'haf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'haf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb0] = (10'hb0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb0] = axis_fifo_inst__DOT__write & (10'hb0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb1] = (10'hb1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb1] = axis_fifo_inst__DOT__write & (10'hb1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb2] = (10'hb2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb2] = axis_fifo_inst__DOT__write & (10'hb2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb3] = (10'hb3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb3] = axis_fifo_inst__DOT__write & (10'hb3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb4] = (10'hb4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb4] = axis_fifo_inst__DOT__write & (10'hb4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb5] = (10'hb5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb5] = axis_fifo_inst__DOT__write & (10'hb5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb6] = (10'hb6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb6] = axis_fifo_inst__DOT__write & (10'hb6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb7] = (10'hb7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb7] = axis_fifo_inst__DOT__write & (10'hb7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb8] = (10'hb8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb8] = axis_fifo_inst__DOT__write & (10'hb8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb9] = (10'hb9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb9] = axis_fifo_inst__DOT__write & (10'hb9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hba] = (10'hba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hba] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hba] = axis_fifo_inst__DOT__write & (10'hba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hba] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hba] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbb] = (10'hbb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbb] = axis_fifo_inst__DOT__write & (10'hbb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbc] = (10'hbc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbc] = axis_fifo_inst__DOT__write & (10'hbc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbd] = (10'hbd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbd] = axis_fifo_inst__DOT__write & (10'hbd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbe] = (10'hbe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbe] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbe] = axis_fifo_inst__DOT__write & (10'hbe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbe] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbe] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbf] = (10'hbf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbf] = axis_fifo_inst__DOT__write & (10'hbf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc0] = (10'hc0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc0] = axis_fifo_inst__DOT__write & (10'hc0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc1] = (10'hc1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc1] = axis_fifo_inst__DOT__write & (10'hc1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc2] = (10'hc2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc2] = axis_fifo_inst__DOT__write & (10'hc2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc3] = (10'hc3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc3] = axis_fifo_inst__DOT__write & (10'hc3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc4] = (10'hc4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc4] = axis_fifo_inst__DOT__write & (10'hc4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc5] = (10'hc5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc5] = axis_fifo_inst__DOT__write & (10'hc5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc6] = (10'hc6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc6] = axis_fifo_inst__DOT__write & (10'hc6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc7] = (10'hc7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc7] = axis_fifo_inst__DOT__write & (10'hc7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc8] = (10'hc8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc8] = axis_fifo_inst__DOT__write & (10'hc8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc9] = (10'hc9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc9] = axis_fifo_inst__DOT__write & (10'hc9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hca] = (10'hca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hca] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hca] = axis_fifo_inst__DOT__write & (10'hca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hca] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hca] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcb] = (10'hcb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcb] = axis_fifo_inst__DOT__write & (10'hcb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcc] = (10'hcc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcc] = axis_fifo_inst__DOT__write & (10'hcc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcd] = (10'hcd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcd] = axis_fifo_inst__DOT__write & (10'hcd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hce] = (10'hce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hce] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hce] = axis_fifo_inst__DOT__write & (10'hce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hce] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hce] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcf] = (10'hcf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcf] = axis_fifo_inst__DOT__write & (10'hcf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd0] = (10'hd0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd0] = axis_fifo_inst__DOT__write & (10'hd0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd1] = (10'hd1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd1] = axis_fifo_inst__DOT__write & (10'hd1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd2] = (10'hd2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd2] = axis_fifo_inst__DOT__write & (10'hd2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd3] = (10'hd3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd3] = axis_fifo_inst__DOT__write & (10'hd3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd4] = (10'hd4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd4] = axis_fifo_inst__DOT__write & (10'hd4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd5] = (10'hd5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd5] = axis_fifo_inst__DOT__write & (10'hd5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd6] = (10'hd6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd6] = axis_fifo_inst__DOT__write & (10'hd6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd7] = (10'hd7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd7] = axis_fifo_inst__DOT__write & (10'hd7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd8] = (10'hd8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd8] = axis_fifo_inst__DOT__write & (10'hd8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd9] = (10'hd9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd9] = axis_fifo_inst__DOT__write & (10'hd9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hda] = (10'hda == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hda] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hda] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hda];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hda] = axis_fifo_inst__DOT__write & (10'hda == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hda] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hda] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hda] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hda];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdb] = (10'hdb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdb] = axis_fifo_inst__DOT__write & (10'hdb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdc] = (10'hdc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdc] = axis_fifo_inst__DOT__write & (10'hdc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdd] = (10'hdd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdd] = axis_fifo_inst__DOT__write & (10'hdd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hde] = (10'hde == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hde] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hde] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hde];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hde] = axis_fifo_inst__DOT__write & (10'hde == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hde] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hde] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hde] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hde];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdf] = (10'hdf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdf] = axis_fifo_inst__DOT__write & (10'hdf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he0] = (10'he0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he0] = axis_fifo_inst__DOT__write & (10'he0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he1] = (10'he1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he1] = axis_fifo_inst__DOT__write & (10'he1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he2] = (10'he2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he2] = axis_fifo_inst__DOT__write & (10'he2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he3] = (10'he3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he3] = axis_fifo_inst__DOT__write & (10'he3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he4] = (10'he4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he4] = axis_fifo_inst__DOT__write & (10'he4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he5] = (10'he5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he5] = axis_fifo_inst__DOT__write & (10'he5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he6] = (10'he6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he6] = axis_fifo_inst__DOT__write & (10'he6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he7] = (10'he7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he7] = axis_fifo_inst__DOT__write & (10'he7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he8] = (10'he8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he8] = axis_fifo_inst__DOT__write & (10'he8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he9] = (10'he9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he9] = axis_fifo_inst__DOT__write & (10'he9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hea] = (10'hea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hea] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hea] = axis_fifo_inst__DOT__write & (10'hea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hea] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hea] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'heb] = (10'heb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'heb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'heb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'heb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'heb] = axis_fifo_inst__DOT__write & (10'heb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'heb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'heb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'heb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'heb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hec] = (10'hec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hec] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hec] = axis_fifo_inst__DOT__write & (10'hec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hec] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hec] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hed] = (10'hed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hed] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hed] = axis_fifo_inst__DOT__write & (10'hed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hed] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hed] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hee] = (10'hee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hee] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hee] = axis_fifo_inst__DOT__write & (10'hee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hee] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hee] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hef] = (10'hef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hef] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hef] = axis_fifo_inst__DOT__write & (10'hef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hef] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hef] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf0] = (10'hf0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf0] = axis_fifo_inst__DOT__write & (10'hf0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf1] = (10'hf1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf1] = axis_fifo_inst__DOT__write & (10'hf1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf2] = (10'hf2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf2] = axis_fifo_inst__DOT__write & (10'hf2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf3] = (10'hf3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf3] = axis_fifo_inst__DOT__write & (10'hf3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf4] = (10'hf4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf4] = axis_fifo_inst__DOT__write & (10'hf4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf5] = (10'hf5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf5] = axis_fifo_inst__DOT__write & (10'hf5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf6] = (10'hf6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf6] = axis_fifo_inst__DOT__write & (10'hf6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf7] = (10'hf7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf7] = axis_fifo_inst__DOT__write & (10'hf7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf8] = (10'hf8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf8] = axis_fifo_inst__DOT__write & (10'hf8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf9] = (10'hf9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf9] = axis_fifo_inst__DOT__write & (10'hf9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfa] = (10'hfa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfa] = axis_fifo_inst__DOT__write & (10'hfa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfb] = (10'hfb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfb] = axis_fifo_inst__DOT__write & (10'hfb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfc] = (10'hfc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfc] = axis_fifo_inst__DOT__write & (10'hfc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfd] = (10'hfd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfd] = axis_fifo_inst__DOT__write & (10'hfd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfe] = (10'hfe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfe] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfe] = axis_fifo_inst__DOT__write & (10'hfe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfe] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfe] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hff] = (10'hff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hff] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hff];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hff] = axis_fifo_inst__DOT__write & (10'hff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hff] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hff] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hff];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h100] = (10'h100 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h100] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h100] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h100];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h100] = axis_fifo_inst__DOT__write & (10'h100 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h100] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h100] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h100] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h100];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h101] = (10'h101 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h101] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h101] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h101];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h101] = axis_fifo_inst__DOT__write & (10'h101 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h101] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h101] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h101] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h101];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h102] = (10'h102 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h102] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h102] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h102];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h102] = axis_fifo_inst__DOT__write & (10'h102 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h102] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h102] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h102] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h102];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h103] = (10'h103 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h103] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h103] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h103];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h103] = axis_fifo_inst__DOT__write & (10'h103 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h103] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h103] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h103] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h103];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h104] = (10'h104 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h104] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h104] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h104];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h104] = axis_fifo_inst__DOT__write & (10'h104 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h104] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h104] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h104] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h104];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h105] = (10'h105 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h105] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h105] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h105];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h105] = axis_fifo_inst__DOT__write & (10'h105 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h105] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h105] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h105] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h105];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h106] = (10'h106 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h106] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h106] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h106];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h106] = axis_fifo_inst__DOT__write & (10'h106 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h106] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h106] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h106] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h106];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h107] = (10'h107 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h107] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h107] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h107];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h107] = axis_fifo_inst__DOT__write & (10'h107 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h107] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h107] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h107] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h107];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h108] = (10'h108 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h108] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h108] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h108];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h108] = axis_fifo_inst__DOT__write & (10'h108 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h108] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h108] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h108] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h108];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h109] = (10'h109 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h109] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h109] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h109];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h109] = axis_fifo_inst__DOT__write & (10'h109 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h109] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h109] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h109] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h109];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10a] = (10'h10a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10a] = axis_fifo_inst__DOT__write & (10'h10a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10b] = (10'h10b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10b] = axis_fifo_inst__DOT__write & (10'h10b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10c] = (10'h10c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10c] = axis_fifo_inst__DOT__write & (10'h10c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10d] = (10'h10d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10d] = axis_fifo_inst__DOT__write & (10'h10d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10e] = (10'h10e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10e] = axis_fifo_inst__DOT__write & (10'h10e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10f] = (10'h10f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10f] = axis_fifo_inst__DOT__write & (10'h10f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h110] = (10'h110 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h110] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h110] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h110];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h110] = axis_fifo_inst__DOT__write & (10'h110 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h110] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h110] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h110] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h110];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h111] = (10'h111 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h111] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h111] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h111];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h111] = axis_fifo_inst__DOT__write & (10'h111 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h111] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h111] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h111] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h111];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h112] = (10'h112 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h112] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h112] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h112];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h112] = axis_fifo_inst__DOT__write & (10'h112 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h112] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h112] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h112] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h112];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h113] = (10'h113 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h113] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h113] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h113];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h113] = axis_fifo_inst__DOT__write & (10'h113 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h113] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h113] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h113] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h113];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h114] = (10'h114 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h114] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h114] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h114];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h114] = axis_fifo_inst__DOT__write & (10'h114 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h114] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h114] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h114] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h114];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h115] = (10'h115 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h115] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h115] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h115];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h115] = axis_fifo_inst__DOT__write & (10'h115 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h115] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h115] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h115] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h115];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h116] = (10'h116 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h116] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h116] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h116];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h116] = axis_fifo_inst__DOT__write & (10'h116 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h116] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h116] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h116] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h116];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h117] = (10'h117 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h117] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h117] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h117];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h117] = axis_fifo_inst__DOT__write & (10'h117 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h117] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h117] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h117] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h117];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h118] = (10'h118 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h118] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h118] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h118];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h118] = axis_fifo_inst__DOT__write & (10'h118 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h118] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h118] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h118] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h118];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h119] = (10'h119 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h119] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h119] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h119];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h119] = axis_fifo_inst__DOT__write & (10'h119 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h119] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h119] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h119] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h119];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11a] = (10'h11a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11a] = axis_fifo_inst__DOT__write & (10'h11a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11b] = (10'h11b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11b] = axis_fifo_inst__DOT__write & (10'h11b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11c] = (10'h11c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11c] = axis_fifo_inst__DOT__write & (10'h11c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11d] = (10'h11d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11d] = axis_fifo_inst__DOT__write & (10'h11d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11e] = (10'h11e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11e] = axis_fifo_inst__DOT__write & (10'h11e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11f] = (10'h11f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11f] = axis_fifo_inst__DOT__write & (10'h11f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h120] = (10'h120 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h120] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h120] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h120];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h120] = axis_fifo_inst__DOT__write & (10'h120 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h120] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h120] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h120] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h120];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h121] = (10'h121 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h121] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h121] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h121];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h121] = axis_fifo_inst__DOT__write & (10'h121 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h121] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h121] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h121] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h121];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h122] = (10'h122 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h122] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h122] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h122];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h122] = axis_fifo_inst__DOT__write & (10'h122 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h122] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h122] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h122] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h122];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h123] = (10'h123 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h123] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h123] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h123];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h123] = axis_fifo_inst__DOT__write & (10'h123 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h123] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h123] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h123] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h123];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h124] = (10'h124 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h124] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h124] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h124];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h124] = axis_fifo_inst__DOT__write & (10'h124 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h124] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h124] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h124] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h124];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h125] = (10'h125 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h125] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h125] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h125];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h125] = axis_fifo_inst__DOT__write & (10'h125 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h125] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h125] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h125] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h125];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h126] = (10'h126 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h126] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h126] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h126];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h126] = axis_fifo_inst__DOT__write & (10'h126 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h126] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h126] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h126] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h126];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h127] = (10'h127 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h127] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h127] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h127];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h127] = axis_fifo_inst__DOT__write & (10'h127 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h127] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h127] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h127] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h127];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h128] = (10'h128 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h128] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h128] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h128];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h128] = axis_fifo_inst__DOT__write & (10'h128 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h128] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h128] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h128] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h128];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h129] = (10'h129 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h129] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h129] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h129];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h129] = axis_fifo_inst__DOT__write & (10'h129 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h129] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h129] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h129] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h129];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12a] = (10'h12a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12a] = axis_fifo_inst__DOT__write & (10'h12a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12b] = (10'h12b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12b] = axis_fifo_inst__DOT__write & (10'h12b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12c] = (10'h12c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12c] = axis_fifo_inst__DOT__write & (10'h12c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12d] = (10'h12d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12d] = axis_fifo_inst__DOT__write & (10'h12d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12e] = (10'h12e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12e] = axis_fifo_inst__DOT__write & (10'h12e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12f] = (10'h12f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12f] = axis_fifo_inst__DOT__write & (10'h12f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h130] = (10'h130 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h130] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h130] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h130];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h130] = axis_fifo_inst__DOT__write & (10'h130 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h130] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h130] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h130] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h130];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h131] = (10'h131 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h131] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h131] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h131];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h131] = axis_fifo_inst__DOT__write & (10'h131 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h131] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h131] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h131] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h131];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h132] = (10'h132 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h132] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h132] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h132];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h132] = axis_fifo_inst__DOT__write & (10'h132 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h132] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h132] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h132] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h132];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h133] = (10'h133 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h133] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h133] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h133];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h133] = axis_fifo_inst__DOT__write & (10'h133 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h133] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h133] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h133] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h133];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h134] = (10'h134 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h134] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h134] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h134];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h134] = axis_fifo_inst__DOT__write & (10'h134 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h134] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h134] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h134] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h134];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h135] = (10'h135 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h135] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h135] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h135];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h135] = axis_fifo_inst__DOT__write & (10'h135 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h135] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h135] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h135] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h135];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h136] = (10'h136 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h136] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h136] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h136];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h136] = axis_fifo_inst__DOT__write & (10'h136 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h136] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h136] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h136] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h136];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h137] = (10'h137 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h137] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h137] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h137];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h137] = axis_fifo_inst__DOT__write & (10'h137 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h137] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h137] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h137] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h137];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h138] = (10'h138 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h138] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h138] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h138];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h138] = axis_fifo_inst__DOT__write & (10'h138 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h138] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h138] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h138] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h138];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h139] = (10'h139 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h139] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h139] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h139];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h139] = axis_fifo_inst__DOT__write & (10'h139 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h139] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h139] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h139] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h139];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13a] = (10'h13a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13a] = axis_fifo_inst__DOT__write & (10'h13a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13b] = (10'h13b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13b] = axis_fifo_inst__DOT__write & (10'h13b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13c] = (10'h13c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13c] = axis_fifo_inst__DOT__write & (10'h13c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13d] = (10'h13d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13d] = axis_fifo_inst__DOT__write & (10'h13d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13e] = (10'h13e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13e] = axis_fifo_inst__DOT__write & (10'h13e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13f] = (10'h13f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13f] = axis_fifo_inst__DOT__write & (10'h13f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h140] = (10'h140 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h140] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h140] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h140];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h140] = axis_fifo_inst__DOT__write & (10'h140 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h140] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h140] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h140] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h140];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h141] = (10'h141 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h141] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h141] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h141];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h141] = axis_fifo_inst__DOT__write & (10'h141 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h141] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h141] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h141] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h141];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h142] = (10'h142 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h142] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h142] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h142];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h142] = axis_fifo_inst__DOT__write & (10'h142 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h142] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h142] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h142] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h142];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h143] = (10'h143 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h143] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h143] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h143];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h143] = axis_fifo_inst__DOT__write & (10'h143 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h143] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h143] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h143] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h143];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h144] = (10'h144 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h144] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h144] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h144];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h144] = axis_fifo_inst__DOT__write & (10'h144 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h144] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h144] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h144] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h144];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h145] = (10'h145 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h145] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h145] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h145];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h145] = axis_fifo_inst__DOT__write & (10'h145 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h145] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h145] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h145] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h145];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h146] = (10'h146 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h146] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h146] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h146];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h146] = axis_fifo_inst__DOT__write & (10'h146 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h146] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h146] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h146] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h146];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h147] = (10'h147 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h147] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h147] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h147];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h147] = axis_fifo_inst__DOT__write & (10'h147 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h147] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h147] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h147] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h147];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h148] = (10'h148 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h148] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h148] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h148];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h148] = axis_fifo_inst__DOT__write & (10'h148 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h148] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h148] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h148] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h148];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h149] = (10'h149 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h149] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h149] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h149];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h149] = axis_fifo_inst__DOT__write & (10'h149 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h149] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h149] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h149] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h149];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14a] = (10'h14a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14a] = axis_fifo_inst__DOT__write & (10'h14a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14b] = (10'h14b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14b] = axis_fifo_inst__DOT__write & (10'h14b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14c] = (10'h14c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14c] = axis_fifo_inst__DOT__write & (10'h14c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14d] = (10'h14d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14d] = axis_fifo_inst__DOT__write & (10'h14d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14e] = (10'h14e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14e] = axis_fifo_inst__DOT__write & (10'h14e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14f] = (10'h14f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14f] = axis_fifo_inst__DOT__write & (10'h14f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h150] = (10'h150 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h150] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h150] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h150];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h150] = axis_fifo_inst__DOT__write & (10'h150 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h150] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h150] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h150] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h150];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h151] = (10'h151 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h151] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h151] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h151];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h151] = axis_fifo_inst__DOT__write & (10'h151 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h151] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h151] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h151] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h151];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h152] = (10'h152 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h152] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h152] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h152];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h152] = axis_fifo_inst__DOT__write & (10'h152 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h152] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h152] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h152] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h152];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h153] = (10'h153 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h153] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h153] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h153];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h153] = axis_fifo_inst__DOT__write & (10'h153 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h153] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h153] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h153] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h153];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h154] = (10'h154 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h154] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h154] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h154];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h154] = axis_fifo_inst__DOT__write & (10'h154 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h154] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h154] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h154] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h154];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h155] = (10'h155 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h155] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h155] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h155];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h155] = axis_fifo_inst__DOT__write & (10'h155 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h155] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h155] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h155] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h155];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h156] = (10'h156 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h156] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h156] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h156];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h156] = axis_fifo_inst__DOT__write & (10'h156 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h156] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h156] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h156] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h156];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h157] = (10'h157 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h157] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h157] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h157];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h157] = axis_fifo_inst__DOT__write & (10'h157 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h157] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h157] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h157] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h157];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h158] = (10'h158 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h158] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h158] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h158];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h158] = axis_fifo_inst__DOT__write & (10'h158 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h158] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h158] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h158] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h158];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h159] = (10'h159 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h159] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h159] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h159];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h159] = axis_fifo_inst__DOT__write & (10'h159 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h159] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h159] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h159] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h159];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15a] = (10'h15a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15a] = axis_fifo_inst__DOT__write & (10'h15a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15b] = (10'h15b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15b] = axis_fifo_inst__DOT__write & (10'h15b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15c] = (10'h15c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15c] = axis_fifo_inst__DOT__write & (10'h15c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15d] = (10'h15d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15d] = axis_fifo_inst__DOT__write & (10'h15d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15e] = (10'h15e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15e] = axis_fifo_inst__DOT__write & (10'h15e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15f] = (10'h15f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15f] = axis_fifo_inst__DOT__write & (10'h15f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h160] = (10'h160 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h160] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h160] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h160];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h160] = axis_fifo_inst__DOT__write & (10'h160 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h160] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h160] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h160] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h160];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h161] = (10'h161 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h161] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h161] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h161];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h161] = axis_fifo_inst__DOT__write & (10'h161 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h161] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h161] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h161] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h161];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h162] = (10'h162 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h162] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h162] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h162];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h162] = axis_fifo_inst__DOT__write & (10'h162 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h162] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h162] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h162] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h162];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h163] = (10'h163 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h163] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h163] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h163];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h163] = axis_fifo_inst__DOT__write & (10'h163 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h163] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h163] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h163] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h163];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h164] = (10'h164 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h164] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h164] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h164];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h164] = axis_fifo_inst__DOT__write & (10'h164 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h164] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h164] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h164] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h164];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h165] = (10'h165 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h165] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h165] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h165];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h165] = axis_fifo_inst__DOT__write & (10'h165 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h165] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h165] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h165] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h165];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h166] = (10'h166 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h166] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h166] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h166];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h166] = axis_fifo_inst__DOT__write & (10'h166 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h166] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h166] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h166] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h166];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h167] = (10'h167 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h167] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h167] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h167];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h167] = axis_fifo_inst__DOT__write & (10'h167 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h167] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h167] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h167] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h167];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h168] = (10'h168 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h168] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h168] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h168];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h168] = axis_fifo_inst__DOT__write & (10'h168 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h168] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h168] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h168] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h168];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h169] = (10'h169 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h169] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h169] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h169];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h169] = axis_fifo_inst__DOT__write & (10'h169 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h169] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h169] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h169] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h169];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16a] = (10'h16a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16a] = axis_fifo_inst__DOT__write & (10'h16a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16b] = (10'h16b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16b] = axis_fifo_inst__DOT__write & (10'h16b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16c] = (10'h16c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16c] = axis_fifo_inst__DOT__write & (10'h16c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16d] = (10'h16d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16d] = axis_fifo_inst__DOT__write & (10'h16d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16e] = (10'h16e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16e] = axis_fifo_inst__DOT__write & (10'h16e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16f] = (10'h16f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16f] = axis_fifo_inst__DOT__write & (10'h16f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h170] = (10'h170 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h170] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h170] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h170];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h170] = axis_fifo_inst__DOT__write & (10'h170 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h170] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h170] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h170] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h170];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h171] = (10'h171 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h171] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h171] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h171];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h171] = axis_fifo_inst__DOT__write & (10'h171 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h171] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h171] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h171] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h171];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h172] = (10'h172 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h172] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h172] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h172];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h172] = axis_fifo_inst__DOT__write & (10'h172 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h172] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h172] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h172] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h172];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h173] = (10'h173 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h173] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h173] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h173];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h173] = axis_fifo_inst__DOT__write & (10'h173 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h173] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h173] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h173] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h173];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h174] = (10'h174 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h174] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h174] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h174];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h174] = axis_fifo_inst__DOT__write & (10'h174 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h174] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h174] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h174] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h174];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h175] = (10'h175 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h175] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h175] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h175];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h175] = axis_fifo_inst__DOT__write & (10'h175 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h175] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h175] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h175] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h175];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h176] = (10'h176 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h176] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h176] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h176];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h176] = axis_fifo_inst__DOT__write & (10'h176 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h176] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h176] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h176] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h176];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h177] = (10'h177 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h177] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h177] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h177];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h177] = axis_fifo_inst__DOT__write & (10'h177 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h177] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h177] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h177] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h177];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h178] = (10'h178 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h178] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h178] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h178];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h178] = axis_fifo_inst__DOT__write & (10'h178 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h178] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h178] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h178] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h178];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h179] = (10'h179 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h179] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h179] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h179];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h179] = axis_fifo_inst__DOT__write & (10'h179 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h179] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h179] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h179] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h179];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17a] = (10'h17a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17a] = axis_fifo_inst__DOT__write & (10'h17a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17b] = (10'h17b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17b] = axis_fifo_inst__DOT__write & (10'h17b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17c] = (10'h17c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17c] = axis_fifo_inst__DOT__write & (10'h17c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17d] = (10'h17d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17d] = axis_fifo_inst__DOT__write & (10'h17d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17e] = (10'h17e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17e] = axis_fifo_inst__DOT__write & (10'h17e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17f] = (10'h17f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17f] = axis_fifo_inst__DOT__write & (10'h17f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h180] = (10'h180 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h180] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h180] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h180];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h180] = axis_fifo_inst__DOT__write & (10'h180 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h180] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h180] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h180] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h180];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h181] = (10'h181 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h181] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h181] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h181];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h181] = axis_fifo_inst__DOT__write & (10'h181 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h181] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h181] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h181] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h181];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h182] = (10'h182 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h182] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h182] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h182];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h182] = axis_fifo_inst__DOT__write & (10'h182 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h182] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h182] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h182] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h182];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h183] = (10'h183 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h183] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h183] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h183];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h183] = axis_fifo_inst__DOT__write & (10'h183 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h183] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h183] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h183] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h183];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h184] = (10'h184 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h184] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h184] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h184];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h184] = axis_fifo_inst__DOT__write & (10'h184 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h184] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h184] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h184] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h184];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h185] = (10'h185 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h185] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h185] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h185];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h185] = axis_fifo_inst__DOT__write & (10'h185 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h185] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h185] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h185] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h185];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h186] = (10'h186 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h186] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h186] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h186];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h186] = axis_fifo_inst__DOT__write & (10'h186 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h186] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h186] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h186] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h186];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h187] = (10'h187 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h187] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h187] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h187];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h187] = axis_fifo_inst__DOT__write & (10'h187 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h187] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h187] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h187] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h187];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h188] = (10'h188 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h188] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h188] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h188];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h188] = axis_fifo_inst__DOT__write & (10'h188 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h188] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h188] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h188] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h188];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h189] = (10'h189 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h189] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h189] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h189];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h189] = axis_fifo_inst__DOT__write & (10'h189 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h189] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h189] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h189] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h189];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18a] = (10'h18a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18a] = axis_fifo_inst__DOT__write & (10'h18a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18b] = (10'h18b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18b] = axis_fifo_inst__DOT__write & (10'h18b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18c] = (10'h18c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18c] = axis_fifo_inst__DOT__write & (10'h18c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18d] = (10'h18d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18d] = axis_fifo_inst__DOT__write & (10'h18d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18e] = (10'h18e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18e] = axis_fifo_inst__DOT__write & (10'h18e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18f] = (10'h18f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18f] = axis_fifo_inst__DOT__write & (10'h18f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h190] = (10'h190 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h190] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h190] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h190];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h190] = axis_fifo_inst__DOT__write & (10'h190 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h190] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h190] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h190] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h190];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h191] = (10'h191 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h191] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h191] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h191];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h191] = axis_fifo_inst__DOT__write & (10'h191 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h191] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h191] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h191] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h191];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h192] = (10'h192 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h192] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h192] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h192];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h192] = axis_fifo_inst__DOT__write & (10'h192 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h192] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h192] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h192] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h192];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h193] = (10'h193 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h193] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h193] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h193];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h193] = axis_fifo_inst__DOT__write & (10'h193 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h193] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h193] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h193] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h193];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h194] = (10'h194 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h194] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h194] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h194];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h194] = axis_fifo_inst__DOT__write & (10'h194 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h194] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h194] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h194] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h194];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h195] = (10'h195 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h195] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h195] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h195];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h195] = axis_fifo_inst__DOT__write & (10'h195 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h195] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h195] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h195] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h195];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h196] = (10'h196 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h196] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h196] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h196];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h196] = axis_fifo_inst__DOT__write & (10'h196 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h196] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h196] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h196] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h196];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h197] = (10'h197 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h197] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h197] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h197];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h197] = axis_fifo_inst__DOT__write & (10'h197 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h197] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h197] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h197] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h197];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h198] = (10'h198 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h198] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h198] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h198];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h198] = axis_fifo_inst__DOT__write & (10'h198 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h198] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h198] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h198] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h198];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h199] = (10'h199 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h199] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h199] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h199];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h199] = axis_fifo_inst__DOT__write & (10'h199 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h199] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h199] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h199] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h199];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19a] = (10'h19a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19a] = axis_fifo_inst__DOT__write & (10'h19a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19b] = (10'h19b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19b] = axis_fifo_inst__DOT__write & (10'h19b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19c] = (10'h19c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19c] = axis_fifo_inst__DOT__write & (10'h19c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19d] = (10'h19d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19d] = axis_fifo_inst__DOT__write & (10'h19d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19e] = (10'h19e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19e] = axis_fifo_inst__DOT__write & (10'h19e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19f] = (10'h19f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19f] = axis_fifo_inst__DOT__write & (10'h19f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a0] = (10'h1a0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a0] = axis_fifo_inst__DOT__write & (10'h1a0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a1] = (10'h1a1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a1] = axis_fifo_inst__DOT__write & (10'h1a1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a2] = (10'h1a2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a2] = axis_fifo_inst__DOT__write & (10'h1a2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a3] = (10'h1a3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a3] = axis_fifo_inst__DOT__write & (10'h1a3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a4] = (10'h1a4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a4] = axis_fifo_inst__DOT__write & (10'h1a4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a5] = (10'h1a5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a5] = axis_fifo_inst__DOT__write & (10'h1a5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a6] = (10'h1a6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a6] = axis_fifo_inst__DOT__write & (10'h1a6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a7] = (10'h1a7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a7] = axis_fifo_inst__DOT__write & (10'h1a7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a8] = (10'h1a8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a8] = axis_fifo_inst__DOT__write & (10'h1a8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a9] = (10'h1a9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a9] = axis_fifo_inst__DOT__write & (10'h1a9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1aa] = (10'h1aa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1aa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1aa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1aa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1aa] = axis_fifo_inst__DOT__write & (10'h1aa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1aa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1aa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1aa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1aa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ab] = (10'h1ab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ab] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ab] = axis_fifo_inst__DOT__write & (10'h1ab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ab] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ab] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ac] = (10'h1ac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ac] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ac] = axis_fifo_inst__DOT__write & (10'h1ac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ac] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ac] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ad] = (10'h1ad == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ad] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ad] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ad];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ad] = axis_fifo_inst__DOT__write & (10'h1ad == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ad] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ad] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ad] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ad];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ae] = (10'h1ae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ae] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ae] = axis_fifo_inst__DOT__write & (10'h1ae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ae] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ae] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1af] = (10'h1af == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1af] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1af] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1af];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1af] = axis_fifo_inst__DOT__write & (10'h1af == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1af] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1af] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1af] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1af];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b0] = (10'h1b0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b0] = axis_fifo_inst__DOT__write & (10'h1b0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b1] = (10'h1b1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b1] = axis_fifo_inst__DOT__write & (10'h1b1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b2] = (10'h1b2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b2] = axis_fifo_inst__DOT__write & (10'h1b2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b3] = (10'h1b3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b3] = axis_fifo_inst__DOT__write & (10'h1b3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b4] = (10'h1b4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b4] = axis_fifo_inst__DOT__write & (10'h1b4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b5] = (10'h1b5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b5] = axis_fifo_inst__DOT__write & (10'h1b5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b6] = (10'h1b6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b6] = axis_fifo_inst__DOT__write & (10'h1b6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b7] = (10'h1b7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b7] = axis_fifo_inst__DOT__write & (10'h1b7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b8] = (10'h1b8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b8] = axis_fifo_inst__DOT__write & (10'h1b8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b9] = (10'h1b9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b9] = axis_fifo_inst__DOT__write & (10'h1b9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ba] = (10'h1ba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ba] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ba] = axis_fifo_inst__DOT__write & (10'h1ba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ba] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ba] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bb] = (10'h1bb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bb] = axis_fifo_inst__DOT__write & (10'h1bb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bc] = (10'h1bc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bc] = axis_fifo_inst__DOT__write & (10'h1bc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bd] = (10'h1bd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bd] = axis_fifo_inst__DOT__write & (10'h1bd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1be] = (10'h1be == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1be] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1be] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1be];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1be] = axis_fifo_inst__DOT__write & (10'h1be == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1be] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1be] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1be] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1be];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bf] = (10'h1bf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bf] = axis_fifo_inst__DOT__write & (10'h1bf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c0] = (10'h1c0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c0] = axis_fifo_inst__DOT__write & (10'h1c0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c1] = (10'h1c1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c1] = axis_fifo_inst__DOT__write & (10'h1c1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c2] = (10'h1c2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c2] = axis_fifo_inst__DOT__write & (10'h1c2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c3] = (10'h1c3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c3] = axis_fifo_inst__DOT__write & (10'h1c3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c4] = (10'h1c4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c4] = axis_fifo_inst__DOT__write & (10'h1c4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c5] = (10'h1c5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c5] = axis_fifo_inst__DOT__write & (10'h1c5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c6] = (10'h1c6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c6] = axis_fifo_inst__DOT__write & (10'h1c6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c7] = (10'h1c7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c7] = axis_fifo_inst__DOT__write & (10'h1c7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c8] = (10'h1c8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c8] = axis_fifo_inst__DOT__write & (10'h1c8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c9] = (10'h1c9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c9] = axis_fifo_inst__DOT__write & (10'h1c9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ca] = (10'h1ca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ca] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ca] = axis_fifo_inst__DOT__write & (10'h1ca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ca] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ca] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cb] = (10'h1cb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cb] = axis_fifo_inst__DOT__write & (10'h1cb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cc] = (10'h1cc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cc] = axis_fifo_inst__DOT__write & (10'h1cc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cd] = (10'h1cd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cd] = axis_fifo_inst__DOT__write & (10'h1cd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ce] = (10'h1ce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ce] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ce] = axis_fifo_inst__DOT__write & (10'h1ce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ce] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ce] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cf] = (10'h1cf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cf] = axis_fifo_inst__DOT__write & (10'h1cf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d0] = (10'h1d0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d0] = axis_fifo_inst__DOT__write & (10'h1d0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d1] = (10'h1d1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d1] = axis_fifo_inst__DOT__write & (10'h1d1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d2] = (10'h1d2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d2] = axis_fifo_inst__DOT__write & (10'h1d2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d3] = (10'h1d3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d3] = axis_fifo_inst__DOT__write & (10'h1d3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d4] = (10'h1d4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d4] = axis_fifo_inst__DOT__write & (10'h1d4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d5] = (10'h1d5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d5] = axis_fifo_inst__DOT__write & (10'h1d5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d6] = (10'h1d6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d6] = axis_fifo_inst__DOT__write & (10'h1d6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d7] = (10'h1d7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d7] = axis_fifo_inst__DOT__write & (10'h1d7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d8] = (10'h1d8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d8] = axis_fifo_inst__DOT__write & (10'h1d8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d9] = (10'h1d9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d9] = axis_fifo_inst__DOT__write & (10'h1d9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1da] = (10'h1da == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1da] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1da] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1da];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1da] = axis_fifo_inst__DOT__write & (10'h1da == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1da] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1da] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1da] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1da];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1db] = (10'h1db == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1db] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1db] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1db];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1db] = axis_fifo_inst__DOT__write & (10'h1db == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1db] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1db] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1db] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1db];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1dc] = (10'h1dc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1dc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1dc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1dc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1dc] = axis_fifo_inst__DOT__write & (10'h1dc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1dc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1dc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1dc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1dc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1dd] = (10'h1dd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1dd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1dd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1dd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1dd] = axis_fifo_inst__DOT__write & (10'h1dd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1dd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1dd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1dd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1dd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1de] = (10'h1de == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1de] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1de] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1de];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1de] = axis_fifo_inst__DOT__write & (10'h1de == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1de] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1de] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1de] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1de];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1df] = (10'h1df == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1df] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1df] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1df];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1df] = axis_fifo_inst__DOT__write & (10'h1df == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1df] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1df] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1df] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1df];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e0] = (10'h1e0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e0] = axis_fifo_inst__DOT__write & (10'h1e0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e1] = (10'h1e1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e1] = axis_fifo_inst__DOT__write & (10'h1e1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e2] = (10'h1e2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e2] = axis_fifo_inst__DOT__write & (10'h1e2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e3] = (10'h1e3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e3] = axis_fifo_inst__DOT__write & (10'h1e3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e4] = (10'h1e4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e4] = axis_fifo_inst__DOT__write & (10'h1e4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e5] = (10'h1e5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e5] = axis_fifo_inst__DOT__write & (10'h1e5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e6] = (10'h1e6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e6] = axis_fifo_inst__DOT__write & (10'h1e6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e7] = (10'h1e7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e7] = axis_fifo_inst__DOT__write & (10'h1e7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e8] = (10'h1e8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e8] = axis_fifo_inst__DOT__write & (10'h1e8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e9] = (10'h1e9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e9] = axis_fifo_inst__DOT__write & (10'h1e9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ea] = (10'h1ea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ea] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ea] = axis_fifo_inst__DOT__write & (10'h1ea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ea] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ea] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1eb] = (10'h1eb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1eb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1eb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1eb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1eb] = axis_fifo_inst__DOT__write & (10'h1eb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1eb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1eb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1eb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1eb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ec] = (10'h1ec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ec] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ec] = axis_fifo_inst__DOT__write & (10'h1ec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ec] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ec] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ed] = (10'h1ed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ed] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ed] = axis_fifo_inst__DOT__write & (10'h1ed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ed] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ed] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ee] = (10'h1ee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ee] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ee] = axis_fifo_inst__DOT__write & (10'h1ee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ee] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ee] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ef] = (10'h1ef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ef] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ef] = axis_fifo_inst__DOT__write & (10'h1ef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ef] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ef] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f0] = (10'h1f0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f0] = axis_fifo_inst__DOT__write & (10'h1f0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f1] = (10'h1f1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f1] = axis_fifo_inst__DOT__write & (10'h1f1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f2] = (10'h1f2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f2] = axis_fifo_inst__DOT__write & (10'h1f2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f3] = (10'h1f3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f3] = axis_fifo_inst__DOT__write & (10'h1f3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f4] = (10'h1f4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f4] = axis_fifo_inst__DOT__write & (10'h1f4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f5] = (10'h1f5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f5] = axis_fifo_inst__DOT__write & (10'h1f5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f6] = (10'h1f6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f6] = axis_fifo_inst__DOT__write & (10'h1f6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f7] = (10'h1f7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f7] = axis_fifo_inst__DOT__write & (10'h1f7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f8] = (10'h1f8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f8] = axis_fifo_inst__DOT__write & (10'h1f8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f9] = (10'h1f9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f9] = axis_fifo_inst__DOT__write & (10'h1f9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fa] = (10'h1fa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fa] = axis_fifo_inst__DOT__write & (10'h1fa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fb] = (10'h1fb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fb] = axis_fifo_inst__DOT__write & (10'h1fb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fc] = (10'h1fc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fc] = axis_fifo_inst__DOT__write & (10'h1fc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fd] = (10'h1fd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fd] = axis_fifo_inst__DOT__write & (10'h1fd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fe] = (10'h1fe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fe] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fe] = axis_fifo_inst__DOT__write & (10'h1fe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fe] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fe] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ff] = (10'h1ff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ff] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ff];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ff] = axis_fifo_inst__DOT__write & (10'h1ff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ff] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ff] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ff];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h200] = (10'h200 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h200] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h200] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h200];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h200] = axis_fifo_inst__DOT__write & (10'h200 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h200] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h200] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h200] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h200];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h201] = (10'h201 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h201] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h201] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h201];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h201] = axis_fifo_inst__DOT__write & (10'h201 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h201] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h201] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h201] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h201];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h202] = (10'h202 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h202] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h202] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h202];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h202] = axis_fifo_inst__DOT__write & (10'h202 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h202] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h202] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h202] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h202];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h203] = (10'h203 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h203] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h203] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h203];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h203] = axis_fifo_inst__DOT__write & (10'h203 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h203] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h203] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h203] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h203];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h204] = (10'h204 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h204] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h204] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h204];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h204] = axis_fifo_inst__DOT__write & (10'h204 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h204] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h204] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h204] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h204];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h205] = (10'h205 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h205] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h205] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h205];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h205] = axis_fifo_inst__DOT__write & (10'h205 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h205] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h205] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h205] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h205];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h206] = (10'h206 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h206] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h206] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h206];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h206] = axis_fifo_inst__DOT__write & (10'h206 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h206] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h206] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h206] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h206];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h207] = (10'h207 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h207] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h207] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h207];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h207] = axis_fifo_inst__DOT__write & (10'h207 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h207] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h207] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h207] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h207];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h208] = (10'h208 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h208] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h208] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h208];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h208] = axis_fifo_inst__DOT__write & (10'h208 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h208] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h208] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h208] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h208];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h209] = (10'h209 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h209] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h209] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h209];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h209] = axis_fifo_inst__DOT__write & (10'h209 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h209] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h209] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h209] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h209];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20a] = (10'h20a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20a] = axis_fifo_inst__DOT__write & (10'h20a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20b] = (10'h20b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20b] = axis_fifo_inst__DOT__write & (10'h20b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20c] = (10'h20c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20c] = axis_fifo_inst__DOT__write & (10'h20c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20d] = (10'h20d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20d] = axis_fifo_inst__DOT__write & (10'h20d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20e] = (10'h20e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20e] = axis_fifo_inst__DOT__write & (10'h20e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20f] = (10'h20f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20f] = axis_fifo_inst__DOT__write & (10'h20f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h210] = (10'h210 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h210] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h210] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h210];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h210] = axis_fifo_inst__DOT__write & (10'h210 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h210] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h210] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h210] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h210];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h211] = (10'h211 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h211] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h211] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h211];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h211] = axis_fifo_inst__DOT__write & (10'h211 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h211] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h211] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h211] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h211];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h212] = (10'h212 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h212] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h212] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h212];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h212] = axis_fifo_inst__DOT__write & (10'h212 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h212] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h212] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h212] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h212];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h213] = (10'h213 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h213] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h213] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h213];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h213] = axis_fifo_inst__DOT__write & (10'h213 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h213] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h213] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h213] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h213];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h214] = (10'h214 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h214] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h214] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h214];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h214] = axis_fifo_inst__DOT__write & (10'h214 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h214] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h214] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h214] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h214];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h215] = (10'h215 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h215] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h215] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h215];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h215] = axis_fifo_inst__DOT__write & (10'h215 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h215] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h215] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h215] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h215];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h216] = (10'h216 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h216] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h216] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h216];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h216] = axis_fifo_inst__DOT__write & (10'h216 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h216] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h216] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h216] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h216];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h217] = (10'h217 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h217] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h217] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h217];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h217] = axis_fifo_inst__DOT__write & (10'h217 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h217] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h217] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h217] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h217];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h218] = (10'h218 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h218] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h218] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h218];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h218] = axis_fifo_inst__DOT__write & (10'h218 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h218] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h218] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h218] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h218];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h219] = (10'h219 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h219] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h219] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h219];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h219] = axis_fifo_inst__DOT__write & (10'h219 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h219] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h219] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h219] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h219];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21a] = (10'h21a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21a] = axis_fifo_inst__DOT__write & (10'h21a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21b] = (10'h21b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21b] = axis_fifo_inst__DOT__write & (10'h21b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21c] = (10'h21c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21c] = axis_fifo_inst__DOT__write & (10'h21c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21d] = (10'h21d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21d] = axis_fifo_inst__DOT__write & (10'h21d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21e] = (10'h21e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21e] = axis_fifo_inst__DOT__write & (10'h21e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21f] = (10'h21f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21f] = axis_fifo_inst__DOT__write & (10'h21f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h220] = (10'h220 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h220] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h220] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h220];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h220] = axis_fifo_inst__DOT__write & (10'h220 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h220] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h220] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h220] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h220];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h221] = (10'h221 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h221] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h221] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h221];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h221] = axis_fifo_inst__DOT__write & (10'h221 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h221] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h221] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h221] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h221];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h222] = (10'h222 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h222] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h222] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h222];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h222] = axis_fifo_inst__DOT__write & (10'h222 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h222] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h222] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h222] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h222];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h223] = (10'h223 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h223] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h223] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h223];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h223] = axis_fifo_inst__DOT__write & (10'h223 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h223] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h223] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h223] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h223];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h224] = (10'h224 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h224] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h224] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h224];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h224] = axis_fifo_inst__DOT__write & (10'h224 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h224] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h224] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h224] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h224];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h225] = (10'h225 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h225] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h225] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h225];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h225] = axis_fifo_inst__DOT__write & (10'h225 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h225] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h225] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h225] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h225];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h226] = (10'h226 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h226] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h226] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h226];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h226] = axis_fifo_inst__DOT__write & (10'h226 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h226] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h226] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h226] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h226];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h227] = (10'h227 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h227] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h227] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h227];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h227] = axis_fifo_inst__DOT__write & (10'h227 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h227] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h227] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h227] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h227];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h228] = (10'h228 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h228] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h228] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h228];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h228] = axis_fifo_inst__DOT__write & (10'h228 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h228] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h228] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h228] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h228];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h229] = (10'h229 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h229] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h229] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h229];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h229] = axis_fifo_inst__DOT__write & (10'h229 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h229] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h229] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h229] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h229];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22a] = (10'h22a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22a] = axis_fifo_inst__DOT__write & (10'h22a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22b] = (10'h22b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22b] = axis_fifo_inst__DOT__write & (10'h22b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22c] = (10'h22c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22c] = axis_fifo_inst__DOT__write & (10'h22c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22d] = (10'h22d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22d] = axis_fifo_inst__DOT__write & (10'h22d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22e] = (10'h22e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22e] = axis_fifo_inst__DOT__write & (10'h22e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22f] = (10'h22f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22f] = axis_fifo_inst__DOT__write & (10'h22f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h230] = (10'h230 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h230] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h230] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h230];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h230] = axis_fifo_inst__DOT__write & (10'h230 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h230] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h230] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h230] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h230];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h231] = (10'h231 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h231] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h231] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h231];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h231] = axis_fifo_inst__DOT__write & (10'h231 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h231] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h231] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h231] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h231];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h232] = (10'h232 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h232] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h232] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h232];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h232] = axis_fifo_inst__DOT__write & (10'h232 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h232] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h232] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h232] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h232];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h233] = (10'h233 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h233] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h233] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h233];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h233] = axis_fifo_inst__DOT__write & (10'h233 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h233] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h233] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h233] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h233];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h234] = (10'h234 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h234] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h234] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h234];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h234] = axis_fifo_inst__DOT__write & (10'h234 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h234] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h234] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h234] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h234];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h235] = (10'h235 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h235] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h235] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h235];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h235] = axis_fifo_inst__DOT__write & (10'h235 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h235] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h235] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h235] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h235];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h236] = (10'h236 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h236] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h236] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h236];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h236] = axis_fifo_inst__DOT__write & (10'h236 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h236] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h236] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h236] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h236];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h237] = (10'h237 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h237] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h237] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h237];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h237] = axis_fifo_inst__DOT__write & (10'h237 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h237] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h237] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h237] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h237];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h238] = (10'h238 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h238] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h238] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h238];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h238] = axis_fifo_inst__DOT__write & (10'h238 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h238] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h238] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h238] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h238];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h239] = (10'h239 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h239] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h239] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h239];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h239] = axis_fifo_inst__DOT__write & (10'h239 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h239] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h239] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h239] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h239];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23a] = (10'h23a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23a] = axis_fifo_inst__DOT__write & (10'h23a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23b] = (10'h23b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23b] = axis_fifo_inst__DOT__write & (10'h23b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23c] = (10'h23c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23c] = axis_fifo_inst__DOT__write & (10'h23c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23d] = (10'h23d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23d] = axis_fifo_inst__DOT__write & (10'h23d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23e] = (10'h23e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23e] = axis_fifo_inst__DOT__write & (10'h23e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23f] = (10'h23f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23f] = axis_fifo_inst__DOT__write & (10'h23f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h240] = (10'h240 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h240] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h240] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h240];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h240] = axis_fifo_inst__DOT__write & (10'h240 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h240] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h240] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h240] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h240];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h241] = (10'h241 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h241] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h241] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h241];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h241] = axis_fifo_inst__DOT__write & (10'h241 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h241] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h241] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h241] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h241];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h242] = (10'h242 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h242] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h242] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h242];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h242] = axis_fifo_inst__DOT__write & (10'h242 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h242] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h242] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h242] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h242];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h243] = (10'h243 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h243] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h243] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h243];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h243] = axis_fifo_inst__DOT__write & (10'h243 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h243] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h243] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h243] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h243];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h244] = (10'h244 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h244] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h244] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h244];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h244] = axis_fifo_inst__DOT__write & (10'h244 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h244] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h244] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h244] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h244];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h245] = (10'h245 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h245] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h245] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h245];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h245] = axis_fifo_inst__DOT__write & (10'h245 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h245] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h245] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h245] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h245];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h246] = (10'h246 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h246] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h246] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h246];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h246] = axis_fifo_inst__DOT__write & (10'h246 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h246] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h246] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h246] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h246];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h247] = (10'h247 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h247] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h247] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h247];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h247] = axis_fifo_inst__DOT__write & (10'h247 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h247] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h247] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h247] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h247];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h248] = (10'h248 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h248] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h248] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h248];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h248] = axis_fifo_inst__DOT__write & (10'h248 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h248] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h248] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h248] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h248];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h249] = (10'h249 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h249] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h249] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h249];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h249] = axis_fifo_inst__DOT__write & (10'h249 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h249] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h249] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h249] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h249];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24a] = (10'h24a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24a] = axis_fifo_inst__DOT__write & (10'h24a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24b] = (10'h24b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24b] = axis_fifo_inst__DOT__write & (10'h24b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24c] = (10'h24c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24c] = axis_fifo_inst__DOT__write & (10'h24c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24d] = (10'h24d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24d] = axis_fifo_inst__DOT__write & (10'h24d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24e] = (10'h24e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24e] = axis_fifo_inst__DOT__write & (10'h24e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24f] = (10'h24f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24f] = axis_fifo_inst__DOT__write & (10'h24f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h250] = (10'h250 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h250] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h250] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h250];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h250] = axis_fifo_inst__DOT__write & (10'h250 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h250] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h250] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h250] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h250];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h251] = (10'h251 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h251] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h251] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h251];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h251] = axis_fifo_inst__DOT__write & (10'h251 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h251] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h251] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h251] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h251];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h252] = (10'h252 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h252] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h252] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h252];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h252] = axis_fifo_inst__DOT__write & (10'h252 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h252] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h252] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h252] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h252];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h253] = (10'h253 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h253] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h253] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h253];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h253] = axis_fifo_inst__DOT__write & (10'h253 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h253] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h253] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h253] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h253];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h254] = (10'h254 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h254] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h254] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h254];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h254] = axis_fifo_inst__DOT__write & (10'h254 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h254] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h254] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h254] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h254];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h255] = (10'h255 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h255] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h255] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h255];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h255] = axis_fifo_inst__DOT__write & (10'h255 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h255] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h255] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h255] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h255];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h256] = (10'h256 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h256] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h256] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h256];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h256] = axis_fifo_inst__DOT__write & (10'h256 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h256] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h256] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h256] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h256];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h257] = (10'h257 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h257] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h257] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h257];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h257] = axis_fifo_inst__DOT__write & (10'h257 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h257] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h257] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h257] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h257];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h258] = (10'h258 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h258] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h258] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h258];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h258] = axis_fifo_inst__DOT__write & (10'h258 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h258] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h258] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h258] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h258];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h259] = (10'h259 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h259] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h259] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h259];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h259] = axis_fifo_inst__DOT__write & (10'h259 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h259] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h259] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h259] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h259];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25a] = (10'h25a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25a] = axis_fifo_inst__DOT__write & (10'h25a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25b] = (10'h25b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25b] = axis_fifo_inst__DOT__write & (10'h25b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25c] = (10'h25c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25c] = axis_fifo_inst__DOT__write & (10'h25c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25d] = (10'h25d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25d] = axis_fifo_inst__DOT__write & (10'h25d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25e] = (10'h25e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25e] = axis_fifo_inst__DOT__write & (10'h25e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25f] = (10'h25f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25f] = axis_fifo_inst__DOT__write & (10'h25f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h260] = (10'h260 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h260] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h260] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h260];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h260] = axis_fifo_inst__DOT__write & (10'h260 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h260] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h260] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h260] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h260];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h261] = (10'h261 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h261] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h261] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h261];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h261] = axis_fifo_inst__DOT__write & (10'h261 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h261] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h261] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h261] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h261];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h262] = (10'h262 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h262] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h262] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h262];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h262] = axis_fifo_inst__DOT__write & (10'h262 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h262] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h262] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h262] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h262];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h263] = (10'h263 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h263] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h263] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h263];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h263] = axis_fifo_inst__DOT__write & (10'h263 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h263] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h263] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h263] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h263];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h264] = (10'h264 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h264] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h264] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h264];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h264] = axis_fifo_inst__DOT__write & (10'h264 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h264] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h264] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h264] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h264];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h265] = (10'h265 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h265] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h265] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h265];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h265] = axis_fifo_inst__DOT__write & (10'h265 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h265] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h265] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h265] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h265];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h266] = (10'h266 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h266] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h266] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h266];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h266] = axis_fifo_inst__DOT__write & (10'h266 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h266] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h266] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h266] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h266];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h267] = (10'h267 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h267] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h267] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h267];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h267] = axis_fifo_inst__DOT__write & (10'h267 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h267] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h267] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h267] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h267];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h268] = (10'h268 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h268] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h268] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h268];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h268] = axis_fifo_inst__DOT__write & (10'h268 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h268] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h268] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h268] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h268];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h269] = (10'h269 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h269] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h269] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h269];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h269] = axis_fifo_inst__DOT__write & (10'h269 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h269] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h269] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h269] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h269];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26a] = (10'h26a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26a] = axis_fifo_inst__DOT__write & (10'h26a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26b] = (10'h26b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26b] = axis_fifo_inst__DOT__write & (10'h26b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26c] = (10'h26c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26c] = axis_fifo_inst__DOT__write & (10'h26c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26d] = (10'h26d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26d] = axis_fifo_inst__DOT__write & (10'h26d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26e] = (10'h26e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26e] = axis_fifo_inst__DOT__write & (10'h26e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26f] = (10'h26f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26f] = axis_fifo_inst__DOT__write & (10'h26f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h270] = (10'h270 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h270] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h270] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h270];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h270] = axis_fifo_inst__DOT__write & (10'h270 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h270] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h270] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h270] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h270];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h271] = (10'h271 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h271] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h271] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h271];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h271] = axis_fifo_inst__DOT__write & (10'h271 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h271] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h271] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h271] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h271];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h272] = (10'h272 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h272] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h272] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h272];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h272] = axis_fifo_inst__DOT__write & (10'h272 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h272] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h272] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h272] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h272];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h273] = (10'h273 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h273] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h273] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h273];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h273] = axis_fifo_inst__DOT__write & (10'h273 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h273] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h273] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h273] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h273];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h274] = (10'h274 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h274] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h274] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h274];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h274] = axis_fifo_inst__DOT__write & (10'h274 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h274] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h274] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h274] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h274];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h275] = (10'h275 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h275] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h275] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h275];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h275] = axis_fifo_inst__DOT__write & (10'h275 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h275] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h275] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h275] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h275];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h276] = (10'h276 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h276] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h276] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h276];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h276] = axis_fifo_inst__DOT__write & (10'h276 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h276] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h276] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h276] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h276];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h277] = (10'h277 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h277] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h277] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h277];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h277] = axis_fifo_inst__DOT__write & (10'h277 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h277] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h277] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h277] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h277];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h278] = (10'h278 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h278] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h278] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h278];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h278] = axis_fifo_inst__DOT__write & (10'h278 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h278] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h278] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h278] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h278];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h279] = (10'h279 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h279] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h279] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h279];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h279] = axis_fifo_inst__DOT__write & (10'h279 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h279] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h279] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h279] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h279];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27a] = (10'h27a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27a] = axis_fifo_inst__DOT__write & (10'h27a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27b] = (10'h27b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27b] = axis_fifo_inst__DOT__write & (10'h27b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27c] = (10'h27c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27c] = axis_fifo_inst__DOT__write & (10'h27c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27d] = (10'h27d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27d] = axis_fifo_inst__DOT__write & (10'h27d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27e] = (10'h27e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27e] = axis_fifo_inst__DOT__write & (10'h27e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27f] = (10'h27f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27f] = axis_fifo_inst__DOT__write & (10'h27f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h280] = (10'h280 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h280] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h280] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h280];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h280] = axis_fifo_inst__DOT__write & (10'h280 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h280] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h280] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h280] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h280];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h281] = (10'h281 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h281] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h281] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h281];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h281] = axis_fifo_inst__DOT__write & (10'h281 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h281] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h281] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h281] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h281];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h282] = (10'h282 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h282] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h282] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h282];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h282] = axis_fifo_inst__DOT__write & (10'h282 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h282] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h282] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h282] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h282];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h283] = (10'h283 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h283] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h283] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h283];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h283] = axis_fifo_inst__DOT__write & (10'h283 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h283] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h283] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h283] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h283];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h284] = (10'h284 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h284] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h284] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h284];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h284] = axis_fifo_inst__DOT__write & (10'h284 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h284] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h284] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h284] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h284];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h285] = (10'h285 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h285] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h285] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h285];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h285] = axis_fifo_inst__DOT__write & (10'h285 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h285] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h285] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h285] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h285];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h286] = (10'h286 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h286] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h286] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h286];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h286] = axis_fifo_inst__DOT__write & (10'h286 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h286] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h286] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h286] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h286];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h287] = (10'h287 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h287] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h287] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h287];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h287] = axis_fifo_inst__DOT__write & (10'h287 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h287] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h287] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h287] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h287];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h288] = (10'h288 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h288] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h288] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h288];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h288] = axis_fifo_inst__DOT__write & (10'h288 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h288] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h288] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h288] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h288];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h289] = (10'h289 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h289] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h289] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h289];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h289] = axis_fifo_inst__DOT__write & (10'h289 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h289] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h289] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h289] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h289];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28a] = (10'h28a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28a] = axis_fifo_inst__DOT__write & (10'h28a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28b] = (10'h28b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28b] = axis_fifo_inst__DOT__write & (10'h28b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28c] = (10'h28c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28c] = axis_fifo_inst__DOT__write & (10'h28c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28d] = (10'h28d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28d] = axis_fifo_inst__DOT__write & (10'h28d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28e] = (10'h28e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28e] = axis_fifo_inst__DOT__write & (10'h28e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28f] = (10'h28f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28f] = axis_fifo_inst__DOT__write & (10'h28f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h290] = (10'h290 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h290] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h290] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h290];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h290] = axis_fifo_inst__DOT__write & (10'h290 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h290] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h290] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h290] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h290];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h291] = (10'h291 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h291] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h291] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h291];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h291] = axis_fifo_inst__DOT__write & (10'h291 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h291] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h291] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h291] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h291];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h292] = (10'h292 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h292] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h292] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h292];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h292] = axis_fifo_inst__DOT__write & (10'h292 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h292] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h292] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h292] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h292];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h293] = (10'h293 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h293] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h293] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h293];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h293] = axis_fifo_inst__DOT__write & (10'h293 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h293] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h293] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h293] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h293];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h294] = (10'h294 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h294] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h294] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h294];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h294] = axis_fifo_inst__DOT__write & (10'h294 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h294] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h294] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h294] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h294];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h295] = (10'h295 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h295] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h295] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h295];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h295] = axis_fifo_inst__DOT__write & (10'h295 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h295] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h295] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h295] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h295];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h296] = (10'h296 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h296] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h296] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h296];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h296] = axis_fifo_inst__DOT__write & (10'h296 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h296] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h296] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h296] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h296];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h297] = (10'h297 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h297] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h297] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h297];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h297] = axis_fifo_inst__DOT__write & (10'h297 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h297] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h297] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h297] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h297];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h298] = (10'h298 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h298] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h298] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h298];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h298] = axis_fifo_inst__DOT__write & (10'h298 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h298] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h298] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h298] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h298];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h299] = (10'h299 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h299] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h299] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h299];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h299] = axis_fifo_inst__DOT__write & (10'h299 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h299] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h299] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h299] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h299];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29a] = (10'h29a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29a] = axis_fifo_inst__DOT__write & (10'h29a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29b] = (10'h29b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29b] = axis_fifo_inst__DOT__write & (10'h29b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29c] = (10'h29c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29c] = axis_fifo_inst__DOT__write & (10'h29c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29d] = (10'h29d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29d] = axis_fifo_inst__DOT__write & (10'h29d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29e] = (10'h29e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29e] = axis_fifo_inst__DOT__write & (10'h29e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29f] = (10'h29f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29f] = axis_fifo_inst__DOT__write & (10'h29f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a0] = (10'h2a0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a0] = axis_fifo_inst__DOT__write & (10'h2a0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a1] = (10'h2a1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a1] = axis_fifo_inst__DOT__write & (10'h2a1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a2] = (10'h2a2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a2] = axis_fifo_inst__DOT__write & (10'h2a2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a3] = (10'h2a3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a3] = axis_fifo_inst__DOT__write & (10'h2a3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a4] = (10'h2a4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a4] = axis_fifo_inst__DOT__write & (10'h2a4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a5] = (10'h2a5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a5] = axis_fifo_inst__DOT__write & (10'h2a5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a6] = (10'h2a6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a6] = axis_fifo_inst__DOT__write & (10'h2a6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a7] = (10'h2a7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a7] = axis_fifo_inst__DOT__write & (10'h2a7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a8] = (10'h2a8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a8] = axis_fifo_inst__DOT__write & (10'h2a8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a9] = (10'h2a9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a9] = axis_fifo_inst__DOT__write & (10'h2a9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2aa] = (10'h2aa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2aa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2aa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2aa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2aa] = axis_fifo_inst__DOT__write & (10'h2aa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2aa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2aa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2aa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2aa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ab] = (10'h2ab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ab] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ab] = axis_fifo_inst__DOT__write & (10'h2ab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ab] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ab] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ac] = (10'h2ac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ac] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ac] = axis_fifo_inst__DOT__write & (10'h2ac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ac] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ac] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ad] = (10'h2ad == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ad] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ad] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ad];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ad] = axis_fifo_inst__DOT__write & (10'h2ad == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ad] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ad] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ad] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ad];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ae] = (10'h2ae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ae] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ae] = axis_fifo_inst__DOT__write & (10'h2ae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ae] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ae] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2af] = (10'h2af == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2af] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2af] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2af];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2af] = axis_fifo_inst__DOT__write & (10'h2af == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2af] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2af] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2af] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2af];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b0] = (10'h2b0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b0] = axis_fifo_inst__DOT__write & (10'h2b0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b1] = (10'h2b1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b1] = axis_fifo_inst__DOT__write & (10'h2b1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b2] = (10'h2b2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b2] = axis_fifo_inst__DOT__write & (10'h2b2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b3] = (10'h2b3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b3] = axis_fifo_inst__DOT__write & (10'h2b3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b4] = (10'h2b4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b4] = axis_fifo_inst__DOT__write & (10'h2b4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b5] = (10'h2b5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b5] = axis_fifo_inst__DOT__write & (10'h2b5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b6] = (10'h2b6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b6] = axis_fifo_inst__DOT__write & (10'h2b6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b7] = (10'h2b7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b7] = axis_fifo_inst__DOT__write & (10'h2b7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b8] = (10'h2b8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b8] = axis_fifo_inst__DOT__write & (10'h2b8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b9] = (10'h2b9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b9] = axis_fifo_inst__DOT__write & (10'h2b9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ba] = (10'h2ba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ba] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ba] = axis_fifo_inst__DOT__write & (10'h2ba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ba] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ba] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bb] = (10'h2bb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bb] = axis_fifo_inst__DOT__write & (10'h2bb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bc] = (10'h2bc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bc] = axis_fifo_inst__DOT__write & (10'h2bc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bd] = (10'h2bd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bd] = axis_fifo_inst__DOT__write & (10'h2bd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2be] = (10'h2be == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2be] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2be] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2be];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2be] = axis_fifo_inst__DOT__write & (10'h2be == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2be] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2be] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2be] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2be];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bf] = (10'h2bf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bf] = axis_fifo_inst__DOT__write & (10'h2bf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c0] = (10'h2c0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c0] = axis_fifo_inst__DOT__write & (10'h2c0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c1] = (10'h2c1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c1] = axis_fifo_inst__DOT__write & (10'h2c1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c2] = (10'h2c2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c2] = axis_fifo_inst__DOT__write & (10'h2c2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c3] = (10'h2c3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c3] = axis_fifo_inst__DOT__write & (10'h2c3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c4] = (10'h2c4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c4] = axis_fifo_inst__DOT__write & (10'h2c4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c5] = (10'h2c5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c5] = axis_fifo_inst__DOT__write & (10'h2c5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c6] = (10'h2c6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c6] = axis_fifo_inst__DOT__write & (10'h2c6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c7] = (10'h2c7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c7] = axis_fifo_inst__DOT__write & (10'h2c7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c8] = (10'h2c8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c8] = axis_fifo_inst__DOT__write & (10'h2c8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c9] = (10'h2c9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c9] = axis_fifo_inst__DOT__write & (10'h2c9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ca] = (10'h2ca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ca] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ca] = axis_fifo_inst__DOT__write & (10'h2ca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ca] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ca] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cb] = (10'h2cb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cb] = axis_fifo_inst__DOT__write & (10'h2cb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cc] = (10'h2cc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cc] = axis_fifo_inst__DOT__write & (10'h2cc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cd] = (10'h2cd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cd] = axis_fifo_inst__DOT__write & (10'h2cd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ce] = (10'h2ce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ce] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ce] = axis_fifo_inst__DOT__write & (10'h2ce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ce] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ce] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cf] = (10'h2cf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cf] = axis_fifo_inst__DOT__write & (10'h2cf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d0] = (10'h2d0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d0] = axis_fifo_inst__DOT__write & (10'h2d0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d1] = (10'h2d1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d1] = axis_fifo_inst__DOT__write & (10'h2d1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d2] = (10'h2d2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d2] = axis_fifo_inst__DOT__write & (10'h2d2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d3] = (10'h2d3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d3] = axis_fifo_inst__DOT__write & (10'h2d3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d4] = (10'h2d4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d4] = axis_fifo_inst__DOT__write & (10'h2d4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d5] = (10'h2d5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d5] = axis_fifo_inst__DOT__write & (10'h2d5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d6] = (10'h2d6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d6] = axis_fifo_inst__DOT__write & (10'h2d6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d7] = (10'h2d7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d7] = axis_fifo_inst__DOT__write & (10'h2d7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d8] = (10'h2d8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d8] = axis_fifo_inst__DOT__write & (10'h2d8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d9] = (10'h2d9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d9] = axis_fifo_inst__DOT__write & (10'h2d9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2da] = (10'h2da == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2da] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2da] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2da];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2da] = axis_fifo_inst__DOT__write & (10'h2da == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2da] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2da] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2da] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2da];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2db] = (10'h2db == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2db] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2db] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2db];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2db] = axis_fifo_inst__DOT__write & (10'h2db == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2db] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2db] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2db] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2db];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2dc] = (10'h2dc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2dc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2dc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2dc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2dc] = axis_fifo_inst__DOT__write & (10'h2dc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2dc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2dc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2dc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2dc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2dd] = (10'h2dd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2dd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2dd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2dd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2dd] = axis_fifo_inst__DOT__write & (10'h2dd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2dd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2dd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2dd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2dd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2de] = (10'h2de == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2de] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2de] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2de];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2de] = axis_fifo_inst__DOT__write & (10'h2de == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2de] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2de] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2de] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2de];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2df] = (10'h2df == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2df] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2df] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2df];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2df] = axis_fifo_inst__DOT__write & (10'h2df == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2df] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2df] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2df] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2df];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e0] = (10'h2e0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e0] = axis_fifo_inst__DOT__write & (10'h2e0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e1] = (10'h2e1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e1] = axis_fifo_inst__DOT__write & (10'h2e1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e2] = (10'h2e2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e2] = axis_fifo_inst__DOT__write & (10'h2e2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e3] = (10'h2e3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e3] = axis_fifo_inst__DOT__write & (10'h2e3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e4] = (10'h2e4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e4] = axis_fifo_inst__DOT__write & (10'h2e4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e5] = (10'h2e5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e5] = axis_fifo_inst__DOT__write & (10'h2e5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e6] = (10'h2e6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e6] = axis_fifo_inst__DOT__write & (10'h2e6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e7] = (10'h2e7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e7] = axis_fifo_inst__DOT__write & (10'h2e7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e8] = (10'h2e8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e8] = axis_fifo_inst__DOT__write & (10'h2e8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e9] = (10'h2e9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e9] = axis_fifo_inst__DOT__write & (10'h2e9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ea] = (10'h2ea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ea] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ea] = axis_fifo_inst__DOT__write & (10'h2ea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ea] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ea] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2eb] = (10'h2eb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2eb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2eb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2eb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2eb] = axis_fifo_inst__DOT__write & (10'h2eb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2eb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2eb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2eb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2eb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ec] = (10'h2ec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ec] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ec] = axis_fifo_inst__DOT__write & (10'h2ec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ec] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ec] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ed] = (10'h2ed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ed] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ed] = axis_fifo_inst__DOT__write & (10'h2ed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ed] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ed] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ee] = (10'h2ee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ee] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ee] = axis_fifo_inst__DOT__write & (10'h2ee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ee] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ee] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ef] = (10'h2ef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ef] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ef] = axis_fifo_inst__DOT__write & (10'h2ef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ef] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ef] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f0] = (10'h2f0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f0] = axis_fifo_inst__DOT__write & (10'h2f0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f1] = (10'h2f1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f1] = axis_fifo_inst__DOT__write & (10'h2f1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f2] = (10'h2f2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f2] = axis_fifo_inst__DOT__write & (10'h2f2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f3] = (10'h2f3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f3] = axis_fifo_inst__DOT__write & (10'h2f3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f4] = (10'h2f4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f4] = axis_fifo_inst__DOT__write & (10'h2f4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f5] = (10'h2f5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f5] = axis_fifo_inst__DOT__write & (10'h2f5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f6] = (10'h2f6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f6] = axis_fifo_inst__DOT__write & (10'h2f6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f7] = (10'h2f7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f7] = axis_fifo_inst__DOT__write & (10'h2f7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f8] = (10'h2f8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f8] = axis_fifo_inst__DOT__write & (10'h2f8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f9] = (10'h2f9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f9] = axis_fifo_inst__DOT__write & (10'h2f9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fa] = (10'h2fa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fa] = axis_fifo_inst__DOT__write & (10'h2fa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fb] = (10'h2fb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fb] = axis_fifo_inst__DOT__write & (10'h2fb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fc] = (10'h2fc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fc] = axis_fifo_inst__DOT__write & (10'h2fc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fd] = (10'h2fd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fd] = axis_fifo_inst__DOT__write & (10'h2fd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fe] = (10'h2fe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fe] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fe] = axis_fifo_inst__DOT__write & (10'h2fe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fe] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fe] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ff] = (10'h2ff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ff] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ff];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ff] = axis_fifo_inst__DOT__write & (10'h2ff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ff] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ff] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ff];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h300] = (10'h300 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h300] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h300] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h300];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h300] = axis_fifo_inst__DOT__write & (10'h300 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h300] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h300] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h300] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h300];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h301] = (10'h301 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h301] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h301] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h301];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h301] = axis_fifo_inst__DOT__write & (10'h301 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h301] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h301] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h301] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h301];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h302] = (10'h302 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h302] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h302] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h302];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h302] = axis_fifo_inst__DOT__write & (10'h302 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h302] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h302] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h302] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h302];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h303] = (10'h303 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h303] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h303] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h303];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h303] = axis_fifo_inst__DOT__write & (10'h303 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h303] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h303] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h303] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h303];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h304] = (10'h304 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h304] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h304] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h304];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h304] = axis_fifo_inst__DOT__write & (10'h304 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h304] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h304] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h304] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h304];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h305] = (10'h305 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h305] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h305] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h305];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h305] = axis_fifo_inst__DOT__write & (10'h305 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h305] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h305] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h305] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h305];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h306] = (10'h306 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h306] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h306] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h306];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h306] = axis_fifo_inst__DOT__write & (10'h306 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h306] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h306] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h306] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h306];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h307] = (10'h307 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h307] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h307] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h307];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h307] = axis_fifo_inst__DOT__write & (10'h307 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h307] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h307] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h307] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h307];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h308] = (10'h308 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h308] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h308] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h308];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h308] = axis_fifo_inst__DOT__write & (10'h308 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h308] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h308] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h308] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h308];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h309] = (10'h309 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h309] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h309] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h309];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h309] = axis_fifo_inst__DOT__write & (10'h309 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h309] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h309] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h309] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h309];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30a] = (10'h30a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30a] = axis_fifo_inst__DOT__write & (10'h30a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30b] = (10'h30b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30b] = axis_fifo_inst__DOT__write & (10'h30b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30c] = (10'h30c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30c] = axis_fifo_inst__DOT__write & (10'h30c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30d] = (10'h30d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30d] = axis_fifo_inst__DOT__write & (10'h30d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30e] = (10'h30e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30e] = axis_fifo_inst__DOT__write & (10'h30e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30f] = (10'h30f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30f] = axis_fifo_inst__DOT__write & (10'h30f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h310] = (10'h310 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h310] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h310] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h310];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h310] = axis_fifo_inst__DOT__write & (10'h310 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h310] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h310] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h310] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h310];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h311] = (10'h311 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h311] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h311] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h311];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h311] = axis_fifo_inst__DOT__write & (10'h311 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h311] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h311] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h311] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h311];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h312] = (10'h312 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h312] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h312] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h312];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h312] = axis_fifo_inst__DOT__write & (10'h312 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h312] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h312] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h312] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h312];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h313] = (10'h313 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h313] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h313] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h313];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h313] = axis_fifo_inst__DOT__write & (10'h313 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h313] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h313] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h313] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h313];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h314] = (10'h314 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h314] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h314] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h314];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h314] = axis_fifo_inst__DOT__write & (10'h314 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h314] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h314] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h314] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h314];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h315] = (10'h315 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h315] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h315] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h315];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h315] = axis_fifo_inst__DOT__write & (10'h315 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h315] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h315] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h315] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h315];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h316] = (10'h316 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h316] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h316] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h316];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h316] = axis_fifo_inst__DOT__write & (10'h316 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h316] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h316] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h316] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h316];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h317] = (10'h317 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h317] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h317] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h317];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h317] = axis_fifo_inst__DOT__write & (10'h317 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h317] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h317] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h317] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h317];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h318] = (10'h318 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h318] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h318] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h318];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h318] = axis_fifo_inst__DOT__write & (10'h318 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h318] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h318] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h318] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h318];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h319] = (10'h319 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h319] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h319] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h319];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h319] = axis_fifo_inst__DOT__write & (10'h319 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h319] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h319] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h319] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h319];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31a] = (10'h31a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31a] = axis_fifo_inst__DOT__write & (10'h31a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31b] = (10'h31b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31b] = axis_fifo_inst__DOT__write & (10'h31b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31c] = (10'h31c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31c] = axis_fifo_inst__DOT__write & (10'h31c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31d] = (10'h31d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31d] = axis_fifo_inst__DOT__write & (10'h31d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31e] = (10'h31e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31e] = axis_fifo_inst__DOT__write & (10'h31e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31f] = (10'h31f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31f] = axis_fifo_inst__DOT__write & (10'h31f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h320] = (10'h320 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h320] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h320] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h320];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h320] = axis_fifo_inst__DOT__write & (10'h320 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h320] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h320] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h320] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h320];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h321] = (10'h321 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h321] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h321] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h321];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h321] = axis_fifo_inst__DOT__write & (10'h321 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h321] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h321] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h321] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h321];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h322] = (10'h322 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h322] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h322] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h322];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h322] = axis_fifo_inst__DOT__write & (10'h322 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h322] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h322] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h322] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h322];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h323] = (10'h323 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h323] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h323] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h323];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h323] = axis_fifo_inst__DOT__write & (10'h323 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h323] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h323] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h323] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h323];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h324] = (10'h324 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h324] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h324] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h324];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h324] = axis_fifo_inst__DOT__write & (10'h324 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h324] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h324] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h324] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h324];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h325] = (10'h325 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h325] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h325] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h325];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h325] = axis_fifo_inst__DOT__write & (10'h325 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h325] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h325] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h325] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h325];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h326] = (10'h326 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h326] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h326] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h326];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h326] = axis_fifo_inst__DOT__write & (10'h326 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h326] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h326] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h326] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h326];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h327] = (10'h327 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h327] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h327] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h327];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h327] = axis_fifo_inst__DOT__write & (10'h327 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h327] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h327] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h327] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h327];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h328] = (10'h328 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h328] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h328] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h328];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h328] = axis_fifo_inst__DOT__write & (10'h328 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h328] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h328] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h328] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h328];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h329] = (10'h329 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h329] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h329] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h329];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h329] = axis_fifo_inst__DOT__write & (10'h329 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h329] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h329] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h329] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h329];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32a] = (10'h32a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32a] = axis_fifo_inst__DOT__write & (10'h32a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32b] = (10'h32b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32b] = axis_fifo_inst__DOT__write & (10'h32b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32c] = (10'h32c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32c] = axis_fifo_inst__DOT__write & (10'h32c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32d] = (10'h32d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32d] = axis_fifo_inst__DOT__write & (10'h32d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32e] = (10'h32e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32e] = axis_fifo_inst__DOT__write & (10'h32e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32f] = (10'h32f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32f] = axis_fifo_inst__DOT__write & (10'h32f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h330] = (10'h330 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h330] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h330] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h330];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h330] = axis_fifo_inst__DOT__write & (10'h330 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h330] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h330] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h330] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h330];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h331] = (10'h331 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h331] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h331] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h331];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h331] = axis_fifo_inst__DOT__write & (10'h331 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h331] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h331] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h331] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h331];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h332] = (10'h332 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h332] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h332] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h332];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h332] = axis_fifo_inst__DOT__write & (10'h332 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h332] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h332] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h332] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h332];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h333] = (10'h333 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h333] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h333] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h333];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h333] = axis_fifo_inst__DOT__write & (10'h333 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h333] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h333] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h333] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h333];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h334] = (10'h334 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h334] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h334] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h334];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h334] = axis_fifo_inst__DOT__write & (10'h334 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h334] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h334] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h334] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h334];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h335] = (10'h335 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h335] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h335] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h335];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h335] = axis_fifo_inst__DOT__write & (10'h335 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h335] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h335] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h335] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h335];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h336] = (10'h336 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h336] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h336] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h336];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h336] = axis_fifo_inst__DOT__write & (10'h336 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h336] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h336] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h336] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h336];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h337] = (10'h337 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h337] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h337] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h337];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h337] = axis_fifo_inst__DOT__write & (10'h337 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h337] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h337] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h337] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h337];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h338] = (10'h338 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h338] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h338] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h338];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h338] = axis_fifo_inst__DOT__write & (10'h338 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h338] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h338] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h338] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h338];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h339] = (10'h339 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h339] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h339] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h339];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h339] = axis_fifo_inst__DOT__write & (10'h339 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h339] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h339] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h339] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h339];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33a] = (10'h33a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33a] = axis_fifo_inst__DOT__write & (10'h33a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33b] = (10'h33b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33b] = axis_fifo_inst__DOT__write & (10'h33b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33c] = (10'h33c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33c] = axis_fifo_inst__DOT__write & (10'h33c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33d] = (10'h33d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33d] = axis_fifo_inst__DOT__write & (10'h33d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33e] = (10'h33e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33e] = axis_fifo_inst__DOT__write & (10'h33e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33f] = (10'h33f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33f] = axis_fifo_inst__DOT__write & (10'h33f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h340] = (10'h340 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h340] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h340] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h340];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h340] = axis_fifo_inst__DOT__write & (10'h340 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h340] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h340] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h340] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h340];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h341] = (10'h341 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h341] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h341] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h341];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h341] = axis_fifo_inst__DOT__write & (10'h341 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h341] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h341] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h341] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h341];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h342] = (10'h342 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h342] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h342] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h342];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h342] = axis_fifo_inst__DOT__write & (10'h342 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h342] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h342] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h342] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h342];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h343] = (10'h343 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h343] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h343] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h343];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h343] = axis_fifo_inst__DOT__write & (10'h343 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h343] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h343] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h343] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h343];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h344] = (10'h344 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h344] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h344] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h344];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h344] = axis_fifo_inst__DOT__write & (10'h344 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h344] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h344] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h344] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h344];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h345] = (10'h345 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h345] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h345] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h345];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h345] = axis_fifo_inst__DOT__write & (10'h345 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h345] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h345] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h345] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h345];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h346] = (10'h346 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h346] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h346] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h346];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h346] = axis_fifo_inst__DOT__write & (10'h346 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h346] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h346] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h346] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h346];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h347] = (10'h347 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h347] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h347] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h347];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h347] = axis_fifo_inst__DOT__write & (10'h347 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h347] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h347] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h347] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h347];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h348] = (10'h348 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h348] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h348] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h348];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h348] = axis_fifo_inst__DOT__write & (10'h348 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h348] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h348] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h348] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h348];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h349] = (10'h349 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h349] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h349] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h349];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h349] = axis_fifo_inst__DOT__write & (10'h349 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h349] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h349] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h349] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h349];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34a] = (10'h34a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34a] = axis_fifo_inst__DOT__write & (10'h34a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34b] = (10'h34b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34b] = axis_fifo_inst__DOT__write & (10'h34b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34c] = (10'h34c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34c] = axis_fifo_inst__DOT__write & (10'h34c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34d] = (10'h34d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34d] = axis_fifo_inst__DOT__write & (10'h34d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34e] = (10'h34e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34e] = axis_fifo_inst__DOT__write & (10'h34e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34f] = (10'h34f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34f] = axis_fifo_inst__DOT__write & (10'h34f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h350] = (10'h350 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h350] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h350] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h350];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h350] = axis_fifo_inst__DOT__write & (10'h350 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h350] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h350] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h350] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h350];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h351] = (10'h351 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h351] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h351] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h351];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h351] = axis_fifo_inst__DOT__write & (10'h351 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h351] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h351] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h351] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h351];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h352] = (10'h352 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h352] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h352] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h352];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h352] = axis_fifo_inst__DOT__write & (10'h352 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h352] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h352] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h352] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h352];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h353] = (10'h353 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h353] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h353] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h353];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h353] = axis_fifo_inst__DOT__write & (10'h353 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h353] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h353] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h353] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h353];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h354] = (10'h354 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h354] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h354] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h354];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h354] = axis_fifo_inst__DOT__write & (10'h354 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h354] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h354] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h354] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h354];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h355] = (10'h355 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h355] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h355] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h355];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h355] = axis_fifo_inst__DOT__write & (10'h355 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h355] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h355] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h355] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h355];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h356] = (10'h356 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h356] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h356] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h356];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h356] = axis_fifo_inst__DOT__write & (10'h356 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h356] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h356] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h356] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h356];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h357] = (10'h357 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h357] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h357] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h357];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h357] = axis_fifo_inst__DOT__write & (10'h357 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h357] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h357] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h357] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h357];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h358] = (10'h358 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h358] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h358] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h358];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h358] = axis_fifo_inst__DOT__write & (10'h358 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h358] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h358] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h358] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h358];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h359] = (10'h359 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h359] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h359] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h359];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h359] = axis_fifo_inst__DOT__write & (10'h359 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h359] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h359] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h359] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h359];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35a] = (10'h35a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35a] = axis_fifo_inst__DOT__write & (10'h35a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35b] = (10'h35b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35b] = axis_fifo_inst__DOT__write & (10'h35b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35c] = (10'h35c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35c] = axis_fifo_inst__DOT__write & (10'h35c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35d] = (10'h35d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35d] = axis_fifo_inst__DOT__write & (10'h35d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35e] = (10'h35e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35e] = axis_fifo_inst__DOT__write & (10'h35e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35f] = (10'h35f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35f] = axis_fifo_inst__DOT__write & (10'h35f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h360] = (10'h360 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h360] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h360] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h360];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h360] = axis_fifo_inst__DOT__write & (10'h360 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h360] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h360] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h360] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h360];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h361] = (10'h361 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h361] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h361] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h361];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h361] = axis_fifo_inst__DOT__write & (10'h361 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h361] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h361] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h361] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h361];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h362] = (10'h362 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h362] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h362] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h362];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h362] = axis_fifo_inst__DOT__write & (10'h362 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h362] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h362] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h362] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h362];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h363] = (10'h363 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h363] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h363] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h363];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h363] = axis_fifo_inst__DOT__write & (10'h363 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h363] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h363] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h363] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h363];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h364] = (10'h364 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h364] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h364] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h364];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h364] = axis_fifo_inst__DOT__write & (10'h364 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h364] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h364] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h364] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h364];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h365] = (10'h365 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h365] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h365] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h365];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h365] = axis_fifo_inst__DOT__write & (10'h365 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h365] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h365] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h365] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h365];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h366] = (10'h366 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h366] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h366] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h366];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h366] = axis_fifo_inst__DOT__write & (10'h366 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h366] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h366] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h366] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h366];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h367] = (10'h367 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h367] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h367] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h367];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h367] = axis_fifo_inst__DOT__write & (10'h367 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h367] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h367] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h367] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h367];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h368] = (10'h368 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h368] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h368] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h368];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h368] = axis_fifo_inst__DOT__write & (10'h368 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h368] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h368] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h368] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h368];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h369] = (10'h369 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h369] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h369] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h369];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h369] = axis_fifo_inst__DOT__write & (10'h369 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h369] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h369] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h369] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h369];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36a] = (10'h36a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36a] = axis_fifo_inst__DOT__write & (10'h36a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36b] = (10'h36b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36b] = axis_fifo_inst__DOT__write & (10'h36b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36c] = (10'h36c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36c] = axis_fifo_inst__DOT__write & (10'h36c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36d] = (10'h36d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36d] = axis_fifo_inst__DOT__write & (10'h36d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36e] = (10'h36e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36e] = axis_fifo_inst__DOT__write & (10'h36e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36f] = (10'h36f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36f] = axis_fifo_inst__DOT__write & (10'h36f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h370] = (10'h370 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h370] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h370] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h370];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h370] = axis_fifo_inst__DOT__write & (10'h370 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h370] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h370] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h370] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h370];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h371] = (10'h371 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h371] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h371] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h371];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h371] = axis_fifo_inst__DOT__write & (10'h371 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h371] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h371] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h371] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h371];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h372] = (10'h372 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h372] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h372] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h372];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h372] = axis_fifo_inst__DOT__write & (10'h372 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h372] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h372] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h372] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h372];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h373] = (10'h373 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h373] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h373] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h373];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h373] = axis_fifo_inst__DOT__write & (10'h373 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h373] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h373] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h373] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h373];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h374] = (10'h374 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h374] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h374] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h374];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h374] = axis_fifo_inst__DOT__write & (10'h374 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h374] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h374] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h374] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h374];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h375] = (10'h375 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h375] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h375] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h375];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h375] = axis_fifo_inst__DOT__write & (10'h375 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h375] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h375] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h375] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h375];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h376] = (10'h376 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h376] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h376] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h376];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h376] = axis_fifo_inst__DOT__write & (10'h376 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h376] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h376] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h376] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h376];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h377] = (10'h377 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h377] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h377] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h377];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h377] = axis_fifo_inst__DOT__write & (10'h377 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h377] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h377] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h377] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h377];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h378] = (10'h378 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h378] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h378] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h378];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h378] = axis_fifo_inst__DOT__write & (10'h378 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h378] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h378] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h378] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h378];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h379] = (10'h379 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h379] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h379] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h379];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h379] = axis_fifo_inst__DOT__write & (10'h379 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h379] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h379] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h379] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h379];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37a] = (10'h37a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37a] = axis_fifo_inst__DOT__write & (10'h37a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37b] = (10'h37b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37b] = axis_fifo_inst__DOT__write & (10'h37b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37c] = (10'h37c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37c] = axis_fifo_inst__DOT__write & (10'h37c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37d] = (10'h37d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37d] = axis_fifo_inst__DOT__write & (10'h37d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37e] = (10'h37e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37e] = axis_fifo_inst__DOT__write & (10'h37e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37f] = (10'h37f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37f] = axis_fifo_inst__DOT__write & (10'h37f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h380] = (10'h380 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h380] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h380] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h380];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h380] = axis_fifo_inst__DOT__write & (10'h380 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h380] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h380] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h380] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h380];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h381] = (10'h381 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h381] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h381] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h381];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h381] = axis_fifo_inst__DOT__write & (10'h381 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h381] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h381] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h381] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h381];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h382] = (10'h382 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h382] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h382] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h382];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h382] = axis_fifo_inst__DOT__write & (10'h382 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h382] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h382] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h382] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h382];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h383] = (10'h383 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h383] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h383] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h383];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h383] = axis_fifo_inst__DOT__write & (10'h383 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h383] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h383] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h383] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h383];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h384] = (10'h384 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h384] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h384] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h384];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h384] = axis_fifo_inst__DOT__write & (10'h384 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h384] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h384] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h384] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h384];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h385] = (10'h385 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h385] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h385] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h385];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h385] = axis_fifo_inst__DOT__write & (10'h385 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h385] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h385] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h385] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h385];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h386] = (10'h386 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h386] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h386] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h386];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h386] = axis_fifo_inst__DOT__write & (10'h386 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h386] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h386] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h386] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h386];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h387] = (10'h387 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h387] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h387] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h387];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h387] = axis_fifo_inst__DOT__write & (10'h387 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h387] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h387] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h387] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h387];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h388] = (10'h388 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h388] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h388] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h388];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h388] = axis_fifo_inst__DOT__write & (10'h388 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h388] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h388] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h388] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h388];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h389] = (10'h389 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h389] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h389] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h389];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h389] = axis_fifo_inst__DOT__write & (10'h389 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h389] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h389] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h389] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h389];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38a] = (10'h38a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38a] = axis_fifo_inst__DOT__write & (10'h38a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38b] = (10'h38b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38b] = axis_fifo_inst__DOT__write & (10'h38b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38c] = (10'h38c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38c] = axis_fifo_inst__DOT__write & (10'h38c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38d] = (10'h38d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38d] = axis_fifo_inst__DOT__write & (10'h38d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38e] = (10'h38e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38e] = axis_fifo_inst__DOT__write & (10'h38e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38f] = (10'h38f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38f] = axis_fifo_inst__DOT__write & (10'h38f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h390] = (10'h390 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h390] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h390] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h390];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h390] = axis_fifo_inst__DOT__write & (10'h390 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h390] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h390] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h390] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h390];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h391] = (10'h391 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h391] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h391] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h391];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h391] = axis_fifo_inst__DOT__write & (10'h391 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h391] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h391] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h391] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h391];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h392] = (10'h392 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h392] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h392] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h392];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h392] = axis_fifo_inst__DOT__write & (10'h392 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h392] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h392] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h392] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h392];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h393] = (10'h393 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h393] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h393] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h393];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h393] = axis_fifo_inst__DOT__write & (10'h393 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h393] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h393] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h393] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h393];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h394] = (10'h394 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h394] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h394] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h394];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h394] = axis_fifo_inst__DOT__write & (10'h394 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h394] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h394] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h394] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h394];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h395] = (10'h395 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h395] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h395] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h395];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h395] = axis_fifo_inst__DOT__write & (10'h395 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h395] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h395] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h395] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h395];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h396] = (10'h396 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h396] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h396] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h396];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h396] = axis_fifo_inst__DOT__write & (10'h396 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h396] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h396] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h396] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h396];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h397] = (10'h397 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h397] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h397] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h397];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h397] = axis_fifo_inst__DOT__write & (10'h397 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h397] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h397] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h397] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h397];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h398] = (10'h398 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h398] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h398] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h398];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h398] = axis_fifo_inst__DOT__write & (10'h398 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h398] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h398] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h398] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h398];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h399] = (10'h399 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h399] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h399] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h399];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h399] = axis_fifo_inst__DOT__write & (10'h399 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h399] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h399] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h399] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h399];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39a] = (10'h39a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39a] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39a] = axis_fifo_inst__DOT__write & (10'h39a == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39a] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39a] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39a] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39a];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39b] = (10'h39b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39b] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39b] = axis_fifo_inst__DOT__write & (10'h39b == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39b] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39b] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39b] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39b];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39c] = (10'h39c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39c] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39c] = axis_fifo_inst__DOT__write & (10'h39c == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39c] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39c] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39c] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39c];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39d] = (10'h39d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39d] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39d] = axis_fifo_inst__DOT__write & (10'h39d == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39d] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39d] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39d] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39d];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39e] = (10'h39e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39e] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39e] = axis_fifo_inst__DOT__write & (10'h39e == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39e] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39e] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39e] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39e];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39f] = (10'h39f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39f] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39f] = axis_fifo_inst__DOT__write & (10'h39f == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39f] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39f] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39f] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39f];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a0] = (10'h3a0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a0] = axis_fifo_inst__DOT__write & (10'h3a0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a1] = (10'h3a1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a1] = axis_fifo_inst__DOT__write & (10'h3a1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a2] = (10'h3a2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a2] = axis_fifo_inst__DOT__write & (10'h3a2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a3] = (10'h3a3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a3] = axis_fifo_inst__DOT__write & (10'h3a3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a4] = (10'h3a4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a4] = axis_fifo_inst__DOT__write & (10'h3a4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a5] = (10'h3a5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a5] = axis_fifo_inst__DOT__write & (10'h3a5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a6] = (10'h3a6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a6] = axis_fifo_inst__DOT__write & (10'h3a6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a7] = (10'h3a7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a7] = axis_fifo_inst__DOT__write & (10'h3a7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a8] = (10'h3a8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a8] = axis_fifo_inst__DOT__write & (10'h3a8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a9] = (10'h3a9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a9] = axis_fifo_inst__DOT__write & (10'h3a9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3aa] = (10'h3aa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3aa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3aa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3aa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3aa] = axis_fifo_inst__DOT__write & (10'h3aa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3aa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3aa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3aa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3aa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ab] = (10'h3ab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ab] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ab] = axis_fifo_inst__DOT__write & (10'h3ab == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ab] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ab] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ab] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ab];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ac] = (10'h3ac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ac] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ac] = axis_fifo_inst__DOT__write & (10'h3ac == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ac] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ac] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ac] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ac];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ad] = (10'h3ad == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ad] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ad] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ad];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ad] = axis_fifo_inst__DOT__write & (10'h3ad == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ad] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ad] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ad] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ad];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ae] = (10'h3ae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ae] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ae] = axis_fifo_inst__DOT__write & (10'h3ae == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ae] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ae] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ae] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ae];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3af] = (10'h3af == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3af] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3af] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3af];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3af] = axis_fifo_inst__DOT__write & (10'h3af == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3af] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3af] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3af] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3af];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b0] = (10'h3b0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b0] = axis_fifo_inst__DOT__write & (10'h3b0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b1] = (10'h3b1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b1] = axis_fifo_inst__DOT__write & (10'h3b1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b2] = (10'h3b2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b2] = axis_fifo_inst__DOT__write & (10'h3b2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b3] = (10'h3b3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b3] = axis_fifo_inst__DOT__write & (10'h3b3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b4] = (10'h3b4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b4] = axis_fifo_inst__DOT__write & (10'h3b4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b5] = (10'h3b5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b5] = axis_fifo_inst__DOT__write & (10'h3b5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b6] = (10'h3b6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b6] = axis_fifo_inst__DOT__write & (10'h3b6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b7] = (10'h3b7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b7] = axis_fifo_inst__DOT__write & (10'h3b7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b8] = (10'h3b8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b8] = axis_fifo_inst__DOT__write & (10'h3b8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b9] = (10'h3b9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b9] = axis_fifo_inst__DOT__write & (10'h3b9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ba] = (10'h3ba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ba] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ba] = axis_fifo_inst__DOT__write & (10'h3ba == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ba] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ba] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ba] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ba];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bb] = (10'h3bb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bb] = axis_fifo_inst__DOT__write & (10'h3bb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bc] = (10'h3bc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bc] = axis_fifo_inst__DOT__write & (10'h3bc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bd] = (10'h3bd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bd] = axis_fifo_inst__DOT__write & (10'h3bd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3be] = (10'h3be == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3be] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3be] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3be];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3be] = axis_fifo_inst__DOT__write & (10'h3be == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3be] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3be] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3be] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3be];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bf] = (10'h3bf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bf] = axis_fifo_inst__DOT__write & (10'h3bf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c0] = (10'h3c0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c0] = axis_fifo_inst__DOT__write & (10'h3c0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c1] = (10'h3c1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c1] = axis_fifo_inst__DOT__write & (10'h3c1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c2] = (10'h3c2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c2] = axis_fifo_inst__DOT__write & (10'h3c2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c3] = (10'h3c3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c3] = axis_fifo_inst__DOT__write & (10'h3c3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c4] = (10'h3c4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c4] = axis_fifo_inst__DOT__write & (10'h3c4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c5] = (10'h3c5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c5] = axis_fifo_inst__DOT__write & (10'h3c5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c6] = (10'h3c6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c6] = axis_fifo_inst__DOT__write & (10'h3c6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c7] = (10'h3c7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c7] = axis_fifo_inst__DOT__write & (10'h3c7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c8] = (10'h3c8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c8] = axis_fifo_inst__DOT__write & (10'h3c8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c9] = (10'h3c9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c9] = axis_fifo_inst__DOT__write & (10'h3c9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ca] = (10'h3ca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ca] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ca] = axis_fifo_inst__DOT__write & (10'h3ca == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ca] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ca] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ca] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ca];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cb] = (10'h3cb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cb] = axis_fifo_inst__DOT__write & (10'h3cb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cc] = (10'h3cc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cc] = axis_fifo_inst__DOT__write & (10'h3cc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cd] = (10'h3cd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cd] = axis_fifo_inst__DOT__write & (10'h3cd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ce] = (10'h3ce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ce] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ce] = axis_fifo_inst__DOT__write & (10'h3ce == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ce] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ce] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ce] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ce];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cf] = (10'h3cf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cf] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cf] = axis_fifo_inst__DOT__write & (10'h3cf == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cf] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cf] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cf] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cf];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d0] = (10'h3d0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d0] = axis_fifo_inst__DOT__write & (10'h3d0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d1] = (10'h3d1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d1] = axis_fifo_inst__DOT__write & (10'h3d1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d2] = (10'h3d2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d2] = axis_fifo_inst__DOT__write & (10'h3d2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d3] = (10'h3d3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d3] = axis_fifo_inst__DOT__write & (10'h3d3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d4] = (10'h3d4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d4] = axis_fifo_inst__DOT__write & (10'h3d4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d5] = (10'h3d5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d5] = axis_fifo_inst__DOT__write & (10'h3d5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d6] = (10'h3d6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d6] = axis_fifo_inst__DOT__write & (10'h3d6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d7] = (10'h3d7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d7] = axis_fifo_inst__DOT__write & (10'h3d7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d8] = (10'h3d8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d8] = axis_fifo_inst__DOT__write & (10'h3d8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d9] = (10'h3d9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d9] = axis_fifo_inst__DOT__write & (10'h3d9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3da] = (10'h3da == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3da] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3da] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3da];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3da] = axis_fifo_inst__DOT__write & (10'h3da == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3da] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3da] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3da] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3da];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3db] = (10'h3db == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3db] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3db] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3db];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3db] = axis_fifo_inst__DOT__write & (10'h3db == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3db] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3db] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3db] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3db];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3dc] = (10'h3dc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3dc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3dc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3dc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3dc] = axis_fifo_inst__DOT__write & (10'h3dc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3dc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3dc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3dc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3dc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3dd] = (10'h3dd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3dd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3dd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3dd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3dd] = axis_fifo_inst__DOT__write & (10'h3dd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3dd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3dd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3dd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3dd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3de] = (10'h3de == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3de] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3de] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3de];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3de] = axis_fifo_inst__DOT__write & (10'h3de == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3de] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3de] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3de] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3de];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3df] = (10'h3df == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3df] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3df] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3df];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3df] = axis_fifo_inst__DOT__write & (10'h3df == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3df] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3df] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3df] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3df];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e0] = (10'h3e0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e0] = axis_fifo_inst__DOT__write & (10'h3e0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e1] = (10'h3e1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e1] = axis_fifo_inst__DOT__write & (10'h3e1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e2] = (10'h3e2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e2] = axis_fifo_inst__DOT__write & (10'h3e2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e3] = (10'h3e3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e3] = axis_fifo_inst__DOT__write & (10'h3e3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e4] = (10'h3e4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e4] = axis_fifo_inst__DOT__write & (10'h3e4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e5] = (10'h3e5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e5] = axis_fifo_inst__DOT__write & (10'h3e5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e6] = (10'h3e6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e6] = axis_fifo_inst__DOT__write & (10'h3e6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e7] = (10'h3e7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e7] = axis_fifo_inst__DOT__write & (10'h3e7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e8] = (10'h3e8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e8] = axis_fifo_inst__DOT__write & (10'h3e8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e9] = (10'h3e9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e9] = axis_fifo_inst__DOT__write & (10'h3e9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ea] = (10'h3ea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ea] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ea] = axis_fifo_inst__DOT__write & (10'h3ea == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ea] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ea] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ea] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ea];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3eb] = (10'h3eb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3eb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3eb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3eb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3eb] = axis_fifo_inst__DOT__write & (10'h3eb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3eb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3eb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3eb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3eb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ec] = (10'h3ec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ec] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ec] = axis_fifo_inst__DOT__write & (10'h3ec == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ec] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ec] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ec] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ec];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ed] = (10'h3ed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ed] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ed] = axis_fifo_inst__DOT__write & (10'h3ed == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ed] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ed] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ed] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ed];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ee] = (10'h3ee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ee] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ee] = axis_fifo_inst__DOT__write & (10'h3ee == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ee] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ee] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ee] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ee];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ef] = (10'h3ef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ef] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ef] = axis_fifo_inst__DOT__write & (10'h3ef == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ef] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ef] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ef] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ef];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f0] = (10'h3f0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f0] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f0] = axis_fifo_inst__DOT__write & (10'h3f0 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f0] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f0] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f0] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f0];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f1] = (10'h3f1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f1] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f1] = axis_fifo_inst__DOT__write & (10'h3f1 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f1] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f1] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f1] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f1];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f2] = (10'h3f2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f2] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f2] = axis_fifo_inst__DOT__write & (10'h3f2 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f2] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f2] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f2] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f2];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f3] = (10'h3f3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f3] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f3] = axis_fifo_inst__DOT__write & (10'h3f3 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f3] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f3] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f3] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f3];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f4] = (10'h3f4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f4] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f4] = axis_fifo_inst__DOT__write & (10'h3f4 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f4] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f4] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f4] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f4];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f5] = (10'h3f5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f5] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f5] = axis_fifo_inst__DOT__write & (10'h3f5 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f5] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f5] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f5] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f5];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f6] = (10'h3f6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f6] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f6] = axis_fifo_inst__DOT__write & (10'h3f6 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f6] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f6] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f6] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f6];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f7] = (10'h3f7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f7] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f7] = axis_fifo_inst__DOT__write & (10'h3f7 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f7] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f7] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f7] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f7];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f8] = (10'h3f8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f8] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f8] = axis_fifo_inst__DOT__write & (10'h3f8 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f8] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f8] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f8] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f8];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f9] = (10'h3f9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f9] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f9] = axis_fifo_inst__DOT__write & (10'h3f9 == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f9] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f9] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f9] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f9];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fa] = (10'h3fa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fa] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fa] = axis_fifo_inst__DOT__write & (10'h3fa == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fa] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fa] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fa] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fa];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fb] = (10'h3fb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fb] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fb] = axis_fifo_inst__DOT__write & (10'h3fb == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fb] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fb] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fb] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fb];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fc] = (10'h3fc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fc] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fc] = axis_fifo_inst__DOT__write & (10'h3fc == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fc] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fc] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fc] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fc];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fd] = (10'h3fd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fd] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fd] = axis_fifo_inst__DOT__write & (10'h3fd == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fd] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fd] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fd] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fd];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fe] = (10'h3fe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fe] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fe] = axis_fifo_inst__DOT__write & (10'h3fe == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fe] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fe] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fe] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fe];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ff] = (10'h3ff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]) & (axis_fifo_inst__DOT__write & axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ff] & ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ff];
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ff] = axis_fifo_inst__DOT__write & (10'h3ff == axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0]);
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ff] = axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ff] | ~axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ff] & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ff];
  assign axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____AV__ = s_axis_tdata__VALID__;
  assign axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____AI__ = axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____ASSIGN__ & ~axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____AV__;
  assign axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____ASSIGN__ = 1'b1;
  assign axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____VALID__ = axis_fifo_inst__DOT__s_axis__BRA__31__03A0__KET____AV__;
  assign axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____PROP__ = 1'b1;
  assign axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____GOOD__ = (rst | axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AI_Q__) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV_Q__) ? (1'b0) : (axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____GOOD_Q__ | axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____PROP_Q__));
  assign axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP__ = axis_fifo_inst__DOT__store_output;
  assign axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD__ = (rst | axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AI_Q__) ? (1'b1) : (
                                                                                (axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV_Q__) ? (1'b0) : (axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD_Q__ | axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP_Q__));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h0] = (10'h0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h0]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1] = (10'h1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2] = (10'h2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3] = (10'h3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4] = (10'h4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5] = (10'h5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6] = (10'h6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7] = (10'h7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8] = (10'h8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9] = (10'h9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha] = (10'ha == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb] = (10'hb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc] = (10'hc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd] = (10'hd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he] = (10'he == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf] = (10'hf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf]) ? (1'b1) : (
                                                                         (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10] = (10'h10 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11] = (10'h11 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12] = (10'h12 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13] = (10'h13 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14] = (10'h14 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15] = (10'h15 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16] = (10'h16 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17] = (10'h17 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18] = (10'h18 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19] = (10'h19 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a] = (10'h1a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b] = (10'h1b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c] = (10'h1c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d] = (10'h1d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e] = (10'h1e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f] = (10'h1f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20] = (10'h20 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21] = (10'h21 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22] = (10'h22 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23] = (10'h23 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24] = (10'h24 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25] = (10'h25 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26] = (10'h26 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27] = (10'h27 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28] = (10'h28 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29] = (10'h29 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a] = (10'h2a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b] = (10'h2b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c] = (10'h2c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d] = (10'h2d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e] = (10'h2e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f] = (10'h2f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30] = (10'h30 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31] = (10'h31 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32] = (10'h32 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33] = (10'h33 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34] = (10'h34 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35] = (10'h35 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36] = (10'h36 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37] = (10'h37 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38] = (10'h38 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39] = (10'h39 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a] = (10'h3a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b] = (10'h3b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c] = (10'h3c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d] = (10'h3d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e] = (10'h3e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f] = (10'h3f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h40] = (10'h40 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h40] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h40]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h40]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h40] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h40]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h41] = (10'h41 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h41] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h41]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h41]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h41] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h41]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h42] = (10'h42 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h42] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h42]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h42]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h42] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h42]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h43] = (10'h43 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h43] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h43]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h43]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h43] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h43]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h44] = (10'h44 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h44] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h44]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h44]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h44] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h44]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h45] = (10'h45 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h45] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h45]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h45]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h45] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h45]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h46] = (10'h46 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h46] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h46]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h46]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h46] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h46]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h47] = (10'h47 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h47] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h47]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h47]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h47] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h47]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h48] = (10'h48 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h48] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h48]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h48]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h48] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h48]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h49] = (10'h49 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h49] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h49]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h49]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h49] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h49]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4a] = (10'h4a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4b] = (10'h4b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4c] = (10'h4c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4d] = (10'h4d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4e] = (10'h4e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4f] = (10'h4f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h50] = (10'h50 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h50] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h50]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h50]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h50] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h50]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h51] = (10'h51 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h51] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h51]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h51]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h51] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h51]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h52] = (10'h52 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h52] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h52]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h52]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h52] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h52]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h53] = (10'h53 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h53] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h53]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h53]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h53] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h53]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h54] = (10'h54 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h54] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h54]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h54]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h54] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h54]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h55] = (10'h55 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h55] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h55]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h55]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h55] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h55]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h56] = (10'h56 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h56] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h56]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h56]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h56] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h56]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h57] = (10'h57 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h57] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h57]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h57]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h57] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h57]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h58] = (10'h58 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h58] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h58]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h58]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h58] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h58]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h59] = (10'h59 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h59] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h59]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h59]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h59] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h59]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5a] = (10'h5a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5b] = (10'h5b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5c] = (10'h5c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5d] = (10'h5d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5e] = (10'h5e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5f] = (10'h5f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h60] = (10'h60 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h60] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h60]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h60]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h60] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h60]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h61] = (10'h61 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h61] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h61]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h61]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h61] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h61]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h62] = (10'h62 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h62] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h62]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h62]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h62] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h62]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h63] = (10'h63 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h63] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h63]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h63]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h63] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h63]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h64] = (10'h64 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h64] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h64]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h64]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h64] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h64]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h65] = (10'h65 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h65] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h65]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h65]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h65] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h65]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h66] = (10'h66 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h66] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h66]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h66]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h66] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h66]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h67] = (10'h67 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h67] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h67]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h67]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h67] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h67]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h68] = (10'h68 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h68] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h68]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h68]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h68] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h68]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h69] = (10'h69 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h69] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h69]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h69]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h69] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h69]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6a] = (10'h6a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6b] = (10'h6b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6c] = (10'h6c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6d] = (10'h6d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6e] = (10'h6e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6f] = (10'h6f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h70] = (10'h70 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h70] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h70]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h70]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h70] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h70]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h71] = (10'h71 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h71] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h71]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h71]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h71] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h71]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h72] = (10'h72 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h72] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h72]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h72]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h72] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h72]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h73] = (10'h73 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h73] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h73]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h73]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h73] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h73]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h74] = (10'h74 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h74] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h74]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h74]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h74] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h74]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h75] = (10'h75 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h75] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h75]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h75]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h75] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h75]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h76] = (10'h76 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h76] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h76]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h76]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h76] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h76]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h77] = (10'h77 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h77] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h77]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h77]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h77] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h77]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h78] = (10'h78 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h78] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h78]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h78]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h78] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h78]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h79] = (10'h79 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h79] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h79]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h79]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h79] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h79]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7a] = (10'h7a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7b] = (10'h7b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7c] = (10'h7c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7d] = (10'h7d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7e] = (10'h7e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7f] = (10'h7f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h80] = (10'h80 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h80] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h80]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h80]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h80] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h80]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h81] = (10'h81 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h81] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h81]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h81]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h81] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h81]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h82] = (10'h82 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h82] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h82]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h82]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h82] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h82]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h83] = (10'h83 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h83] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h83]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h83]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h83] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h83]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h84] = (10'h84 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h84] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h84]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h84]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h84] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h84]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h85] = (10'h85 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h85] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h85]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h85]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h85] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h85]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h86] = (10'h86 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h86] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h86]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h86]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h86] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h86]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h87] = (10'h87 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h87] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h87]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h87]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h87] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h87]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h88] = (10'h88 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h88] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h88]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h88]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h88] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h88]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h89] = (10'h89 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h89] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h89]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h89]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h89] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h89]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8a] = (10'h8a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8b] = (10'h8b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8c] = (10'h8c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8d] = (10'h8d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8e] = (10'h8e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8f] = (10'h8f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h90] = (10'h90 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h90] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h90]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h90]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h90] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h90]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h91] = (10'h91 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h91] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h91]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h91]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h91] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h91]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h92] = (10'h92 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h92] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h92]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h92]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h92] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h92]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h93] = (10'h93 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h93] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h93]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h93]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h93] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h93]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h94] = (10'h94 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h94] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h94]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h94]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h94] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h94]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h95] = (10'h95 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h95] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h95]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h95]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h95] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h95]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h96] = (10'h96 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h96] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h96]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h96]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h96] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h96]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h97] = (10'h97 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h97] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h97]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h97]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h97] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h97]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h98] = (10'h98 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h98] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h98]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h98]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h98] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h98]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h99] = (10'h99 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h99] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h99]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h99]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h99] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h99]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9a] = (10'h9a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9a]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9b] = (10'h9b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9b]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9c] = (10'h9c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9c]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9d] = (10'h9d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9d]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9e] = (10'h9e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9e]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9f] = (10'h9f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9f]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha0] = (10'ha0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha0]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha1] = (10'ha1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha1]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha2] = (10'ha2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha2]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha3] = (10'ha3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha3]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha4] = (10'ha4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha4]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha5] = (10'ha5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha5]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha6] = (10'ha6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha6]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha7] = (10'ha7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha7]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha8] = (10'ha8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha8]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha9] = (10'ha9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha9]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'haa] = (10'haa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'haa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'haa]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'haa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'haa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'haa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hab] = (10'hab == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hab] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hab]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hab]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hab] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hab]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hac] = (10'hac == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hac] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hac]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hac]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hac] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hac]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'had] = (10'had == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'had] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'had]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'had]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'had] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'had]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hae] = (10'hae == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hae] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hae]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hae]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hae] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hae]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'haf] = (10'haf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'haf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'haf]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'haf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'haf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'haf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb0] = (10'hb0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb0]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb1] = (10'hb1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb1]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb2] = (10'hb2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb2]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb3] = (10'hb3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb3]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb4] = (10'hb4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb4]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb5] = (10'hb5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb5]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb6] = (10'hb6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb6]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb7] = (10'hb7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb7]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb8] = (10'hb8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb8]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb9] = (10'hb9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb9]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hba] = (10'hba == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hba] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hba]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hba]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hba] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hba]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbb] = (10'hbb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbb]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbc] = (10'hbc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbc]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbd] = (10'hbd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbd]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbe] = (10'hbe == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbe] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbe]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbe]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbe] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbe]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbf] = (10'hbf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbf]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc0] = (10'hc0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc0]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc1] = (10'hc1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc1]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc2] = (10'hc2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc2]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc3] = (10'hc3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc3]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc4] = (10'hc4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc4]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc5] = (10'hc5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc5]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc6] = (10'hc6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc6]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc7] = (10'hc7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc7]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc8] = (10'hc8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc8]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc9] = (10'hc9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc9]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hca] = (10'hca == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hca] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hca]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hca]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hca] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hca]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcb] = (10'hcb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcb]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcc] = (10'hcc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcc]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcd] = (10'hcd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcd]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hce] = (10'hce == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hce] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hce]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hce]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hce] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hce]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcf] = (10'hcf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcf]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd0] = (10'hd0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd0]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd1] = (10'hd1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd1]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd2] = (10'hd2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd2]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd3] = (10'hd3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd3]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd4] = (10'hd4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd4]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd5] = (10'hd5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd5]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd6] = (10'hd6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd6]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd7] = (10'hd7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd7]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd8] = (10'hd8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd8]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd9] = (10'hd9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd9]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hda] = (10'hda == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hda] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hda]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hda]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hda] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hda]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdb] = (10'hdb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdb]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdc] = (10'hdc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdc]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdd] = (10'hdd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdd]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hde] = (10'hde == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hde] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hde]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hde]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hde] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hde]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdf] = (10'hdf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdf]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he0] = (10'he0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he0]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he1] = (10'he1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he1]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he2] = (10'he2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he2]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he3] = (10'he3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he3]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he4] = (10'he4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he4]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he5] = (10'he5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he5]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he6] = (10'he6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he6]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he7] = (10'he7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he7]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he8] = (10'he8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he8]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he9] = (10'he9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he9]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hea] = (10'hea == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hea] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hea]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hea]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hea] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hea]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'heb] = (10'heb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'heb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'heb]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'heb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'heb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'heb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hec] = (10'hec == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hec] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hec]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hec]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hec] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hec]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hed] = (10'hed == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hed] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hed]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hed]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hed] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hed]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hee] = (10'hee == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hee] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hee]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hee]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hee] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hee]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hef] = (10'hef == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hef] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hef]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hef]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hef] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hef]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf0] = (10'hf0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf0]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf1] = (10'hf1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf1]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf2] = (10'hf2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf2]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf3] = (10'hf3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf3]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf4] = (10'hf4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf4]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf5] = (10'hf5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf5]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf6] = (10'hf6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf6]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf7] = (10'hf7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf7]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf8] = (10'hf8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf8]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf9] = (10'hf9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf9]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfa] = (10'hfa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfa]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfb] = (10'hfb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfb]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfc] = (10'hfc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfc]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfd] = (10'hfd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfd]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfe] = (10'hfe == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfe] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfe]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfe]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfe] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfe]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hff] = (10'hff == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hff] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hff]) ? (1'b1) : (
                                                                          (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hff]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hff] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hff]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h100] = (10'h100 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h100] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h100]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h100]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h100] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h100]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h101] = (10'h101 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h101] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h101]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h101]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h101] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h101]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h102] = (10'h102 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h102] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h102]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h102]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h102] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h102]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h103] = (10'h103 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h103] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h103]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h103]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h103] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h103]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h104] = (10'h104 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h104] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h104]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h104]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h104] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h104]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h105] = (10'h105 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h105] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h105]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h105]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h105] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h105]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h106] = (10'h106 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h106] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h106]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h106]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h106] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h106]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h107] = (10'h107 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h107] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h107]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h107]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h107] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h107]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h108] = (10'h108 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h108] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h108]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h108]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h108] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h108]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h109] = (10'h109 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h109] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h109]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h109]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h109] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h109]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10a] = (10'h10a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10b] = (10'h10b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10c] = (10'h10c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10d] = (10'h10d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10e] = (10'h10e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10f] = (10'h10f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h110] = (10'h110 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h110] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h110]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h110]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h110] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h110]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h111] = (10'h111 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h111] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h111]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h111]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h111] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h111]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h112] = (10'h112 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h112] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h112]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h112]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h112] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h112]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h113] = (10'h113 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h113] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h113]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h113]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h113] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h113]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h114] = (10'h114 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h114] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h114]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h114]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h114] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h114]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h115] = (10'h115 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h115] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h115]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h115]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h115] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h115]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h116] = (10'h116 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h116] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h116]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h116]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h116] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h116]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h117] = (10'h117 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h117] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h117]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h117]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h117] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h117]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h118] = (10'h118 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h118] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h118]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h118]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h118] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h118]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h119] = (10'h119 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h119] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h119]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h119]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h119] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h119]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11a] = (10'h11a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11b] = (10'h11b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11c] = (10'h11c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11d] = (10'h11d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11e] = (10'h11e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11f] = (10'h11f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h120] = (10'h120 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h120] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h120]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h120]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h120] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h120]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h121] = (10'h121 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h121] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h121]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h121]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h121] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h121]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h122] = (10'h122 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h122] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h122]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h122]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h122] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h122]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h123] = (10'h123 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h123] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h123]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h123]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h123] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h123]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h124] = (10'h124 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h124] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h124]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h124]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h124] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h124]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h125] = (10'h125 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h125] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h125]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h125]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h125] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h125]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h126] = (10'h126 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h126] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h126]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h126]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h126] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h126]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h127] = (10'h127 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h127] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h127]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h127]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h127] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h127]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h128] = (10'h128 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h128] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h128]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h128]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h128] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h128]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h129] = (10'h129 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h129] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h129]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h129]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h129] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h129]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12a] = (10'h12a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12b] = (10'h12b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12c] = (10'h12c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12d] = (10'h12d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12e] = (10'h12e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12f] = (10'h12f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h130] = (10'h130 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h130] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h130]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h130]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h130] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h130]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h131] = (10'h131 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h131] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h131]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h131]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h131] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h131]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h132] = (10'h132 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h132] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h132]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h132]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h132] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h132]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h133] = (10'h133 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h133] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h133]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h133]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h133] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h133]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h134] = (10'h134 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h134] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h134]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h134]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h134] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h134]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h135] = (10'h135 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h135] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h135]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h135]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h135] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h135]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h136] = (10'h136 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h136] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h136]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h136]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h136] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h136]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h137] = (10'h137 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h137] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h137]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h137]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h137] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h137]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h138] = (10'h138 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h138] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h138]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h138]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h138] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h138]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h139] = (10'h139 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h139] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h139]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h139]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h139] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h139]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13a] = (10'h13a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13b] = (10'h13b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13c] = (10'h13c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13d] = (10'h13d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13e] = (10'h13e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13f] = (10'h13f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h140] = (10'h140 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h140] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h140]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h140]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h140] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h140]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h141] = (10'h141 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h141] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h141]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h141]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h141] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h141]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h142] = (10'h142 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h142] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h142]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h142]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h142] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h142]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h143] = (10'h143 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h143] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h143]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h143]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h143] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h143]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h144] = (10'h144 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h144] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h144]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h144]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h144] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h144]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h145] = (10'h145 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h145] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h145]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h145]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h145] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h145]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h146] = (10'h146 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h146] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h146]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h146]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h146] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h146]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h147] = (10'h147 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h147] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h147]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h147]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h147] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h147]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h148] = (10'h148 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h148] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h148]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h148]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h148] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h148]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h149] = (10'h149 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h149] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h149]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h149]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h149] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h149]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14a] = (10'h14a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14b] = (10'h14b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14c] = (10'h14c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14d] = (10'h14d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14e] = (10'h14e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14f] = (10'h14f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h150] = (10'h150 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h150] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h150]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h150]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h150] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h150]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h151] = (10'h151 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h151] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h151]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h151]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h151] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h151]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h152] = (10'h152 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h152] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h152]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h152]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h152] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h152]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h153] = (10'h153 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h153] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h153]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h153]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h153] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h153]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h154] = (10'h154 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h154] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h154]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h154]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h154] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h154]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h155] = (10'h155 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h155] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h155]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h155]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h155] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h155]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h156] = (10'h156 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h156] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h156]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h156]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h156] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h156]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h157] = (10'h157 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h157] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h157]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h157]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h157] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h157]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h158] = (10'h158 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h158] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h158]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h158]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h158] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h158]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h159] = (10'h159 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h159] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h159]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h159]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h159] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h159]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15a] = (10'h15a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15b] = (10'h15b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15c] = (10'h15c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15d] = (10'h15d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15e] = (10'h15e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15f] = (10'h15f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h160] = (10'h160 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h160] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h160]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h160]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h160] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h160]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h161] = (10'h161 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h161] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h161]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h161]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h161] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h161]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h162] = (10'h162 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h162] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h162]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h162]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h162] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h162]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h163] = (10'h163 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h163] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h163]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h163]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h163] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h163]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h164] = (10'h164 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h164] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h164]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h164]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h164] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h164]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h165] = (10'h165 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h165] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h165]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h165]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h165] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h165]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h166] = (10'h166 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h166] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h166]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h166]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h166] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h166]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h167] = (10'h167 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h167] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h167]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h167]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h167] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h167]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h168] = (10'h168 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h168] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h168]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h168]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h168] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h168]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h169] = (10'h169 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h169] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h169]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h169]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h169] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h169]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16a] = (10'h16a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16b] = (10'h16b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16c] = (10'h16c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16d] = (10'h16d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16e] = (10'h16e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16f] = (10'h16f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h170] = (10'h170 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h170] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h170]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h170]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h170] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h170]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h171] = (10'h171 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h171] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h171]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h171]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h171] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h171]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h172] = (10'h172 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h172] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h172]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h172]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h172] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h172]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h173] = (10'h173 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h173] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h173]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h173]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h173] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h173]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h174] = (10'h174 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h174] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h174]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h174]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h174] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h174]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h175] = (10'h175 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h175] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h175]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h175]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h175] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h175]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h176] = (10'h176 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h176] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h176]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h176]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h176] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h176]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h177] = (10'h177 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h177] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h177]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h177]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h177] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h177]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h178] = (10'h178 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h178] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h178]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h178]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h178] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h178]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h179] = (10'h179 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h179] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h179]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h179]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h179] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h179]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17a] = (10'h17a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17b] = (10'h17b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17c] = (10'h17c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17d] = (10'h17d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17e] = (10'h17e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17f] = (10'h17f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h180] = (10'h180 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h180] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h180]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h180]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h180] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h180]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h181] = (10'h181 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h181] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h181]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h181]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h181] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h181]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h182] = (10'h182 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h182] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h182]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h182]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h182] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h182]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h183] = (10'h183 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h183] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h183]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h183]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h183] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h183]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h184] = (10'h184 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h184] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h184]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h184]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h184] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h184]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h185] = (10'h185 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h185] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h185]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h185]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h185] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h185]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h186] = (10'h186 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h186] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h186]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h186]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h186] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h186]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h187] = (10'h187 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h187] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h187]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h187]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h187] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h187]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h188] = (10'h188 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h188] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h188]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h188]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h188] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h188]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h189] = (10'h189 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h189] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h189]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h189]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h189] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h189]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18a] = (10'h18a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18b] = (10'h18b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18c] = (10'h18c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18d] = (10'h18d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18e] = (10'h18e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18f] = (10'h18f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h190] = (10'h190 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h190] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h190]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h190]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h190] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h190]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h191] = (10'h191 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h191] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h191]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h191]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h191] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h191]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h192] = (10'h192 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h192] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h192]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h192]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h192] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h192]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h193] = (10'h193 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h193] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h193]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h193]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h193] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h193]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h194] = (10'h194 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h194] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h194]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h194]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h194] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h194]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h195] = (10'h195 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h195] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h195]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h195]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h195] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h195]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h196] = (10'h196 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h196] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h196]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h196]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h196] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h196]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h197] = (10'h197 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h197] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h197]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h197]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h197] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h197]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h198] = (10'h198 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h198] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h198]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h198]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h198] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h198]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h199] = (10'h199 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h199] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h199]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h199]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h199] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h199]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19a] = (10'h19a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19b] = (10'h19b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19c] = (10'h19c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19d] = (10'h19d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19e] = (10'h19e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19f] = (10'h19f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a0] = (10'h1a0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a1] = (10'h1a1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a2] = (10'h1a2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a3] = (10'h1a3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a4] = (10'h1a4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a5] = (10'h1a5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a6] = (10'h1a6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a7] = (10'h1a7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a8] = (10'h1a8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a9] = (10'h1a9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1aa] = (10'h1aa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1aa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1aa]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1aa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1aa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1aa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ab] = (10'h1ab == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ab] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ab]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ab]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ab] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ab]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ac] = (10'h1ac == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ac] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ac]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ac]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ac] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ac]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ad] = (10'h1ad == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ad] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ad]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ad]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ad] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ad]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ae] = (10'h1ae == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ae] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ae]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ae]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ae] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ae]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1af] = (10'h1af == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1af] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1af]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1af]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1af] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1af]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b0] = (10'h1b0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b1] = (10'h1b1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b2] = (10'h1b2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b3] = (10'h1b3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b4] = (10'h1b4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b5] = (10'h1b5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b6] = (10'h1b6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b7] = (10'h1b7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b8] = (10'h1b8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b9] = (10'h1b9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ba] = (10'h1ba == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ba] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ba]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ba]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ba] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ba]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bb] = (10'h1bb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bc] = (10'h1bc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bd] = (10'h1bd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1be] = (10'h1be == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1be] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1be]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1be]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1be] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1be]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bf] = (10'h1bf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bf]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c0] = (10'h1c0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c1] = (10'h1c1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c2] = (10'h1c2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c3] = (10'h1c3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c4] = (10'h1c4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c5] = (10'h1c5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c6] = (10'h1c6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c7] = (10'h1c7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c8] = (10'h1c8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c9] = (10'h1c9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ca] = (10'h1ca == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ca] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ca]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ca]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ca] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ca]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cb] = (10'h1cb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cc] = (10'h1cc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cd] = (10'h1cd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ce] = (10'h1ce == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ce] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ce]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ce]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ce] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ce]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cf] = (10'h1cf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cf]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d0] = (10'h1d0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d1] = (10'h1d1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d2] = (10'h1d2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d3] = (10'h1d3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d4] = (10'h1d4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d5] = (10'h1d5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d6] = (10'h1d6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d7] = (10'h1d7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d8] = (10'h1d8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d9] = (10'h1d9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1da] = (10'h1da == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1da] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1da]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1da]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1da] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1da]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1db] = (10'h1db == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1db] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1db]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1db]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1db] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1db]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1dc] = (10'h1dc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1dc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1dc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1dc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1dc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1dc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1dd] = (10'h1dd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1dd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1dd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1dd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1dd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1dd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1de] = (10'h1de == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1de] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1de]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1de]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1de] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1de]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1df] = (10'h1df == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1df] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1df]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1df]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1df] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1df]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e0] = (10'h1e0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e1] = (10'h1e1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e2] = (10'h1e2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e3] = (10'h1e3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e4] = (10'h1e4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e5] = (10'h1e5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e6] = (10'h1e6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e7] = (10'h1e7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e8] = (10'h1e8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e9] = (10'h1e9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ea] = (10'h1ea == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ea] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ea]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ea]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ea] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ea]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1eb] = (10'h1eb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1eb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1eb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1eb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1eb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1eb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ec] = (10'h1ec == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ec] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ec]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ec]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ec] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ec]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ed] = (10'h1ed == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ed] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ed]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ed]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ed] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ed]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ee] = (10'h1ee == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ee] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ee]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ee]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ee] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ee]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ef] = (10'h1ef == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ef] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ef]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ef]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ef] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ef]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f0] = (10'h1f0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f1] = (10'h1f1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f2] = (10'h1f2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f3] = (10'h1f3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f4] = (10'h1f4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f5] = (10'h1f5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f6] = (10'h1f6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f7] = (10'h1f7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f8] = (10'h1f8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f9] = (10'h1f9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fa] = (10'h1fa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fa]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fb] = (10'h1fb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fc] = (10'h1fc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fd] = (10'h1fd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fe] = (10'h1fe == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fe] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fe]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fe]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fe] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fe]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ff] = (10'h1ff == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ff] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ff]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ff]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ff] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ff]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h200] = (10'h200 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h200] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h200]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h200]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h200] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h200]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h201] = (10'h201 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h201] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h201]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h201]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h201] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h201]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h202] = (10'h202 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h202] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h202]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h202]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h202] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h202]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h203] = (10'h203 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h203] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h203]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h203]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h203] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h203]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h204] = (10'h204 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h204] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h204]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h204]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h204] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h204]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h205] = (10'h205 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h205] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h205]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h205]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h205] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h205]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h206] = (10'h206 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h206] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h206]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h206]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h206] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h206]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h207] = (10'h207 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h207] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h207]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h207]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h207] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h207]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h208] = (10'h208 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h208] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h208]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h208]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h208] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h208]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h209] = (10'h209 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h209] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h209]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h209]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h209] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h209]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20a] = (10'h20a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20b] = (10'h20b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20c] = (10'h20c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20d] = (10'h20d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20e] = (10'h20e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20f] = (10'h20f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h210] = (10'h210 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h210] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h210]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h210]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h210] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h210]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h211] = (10'h211 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h211] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h211]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h211]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h211] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h211]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h212] = (10'h212 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h212] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h212]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h212]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h212] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h212]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h213] = (10'h213 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h213] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h213]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h213]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h213] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h213]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h214] = (10'h214 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h214] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h214]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h214]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h214] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h214]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h215] = (10'h215 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h215] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h215]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h215]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h215] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h215]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h216] = (10'h216 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h216] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h216]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h216]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h216] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h216]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h217] = (10'h217 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h217] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h217]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h217]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h217] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h217]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h218] = (10'h218 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h218] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h218]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h218]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h218] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h218]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h219] = (10'h219 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h219] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h219]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h219]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h219] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h219]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21a] = (10'h21a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21b] = (10'h21b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21c] = (10'h21c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21d] = (10'h21d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21e] = (10'h21e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21f] = (10'h21f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h220] = (10'h220 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h220] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h220]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h220]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h220] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h220]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h221] = (10'h221 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h221] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h221]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h221]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h221] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h221]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h222] = (10'h222 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h222] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h222]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h222]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h222] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h222]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h223] = (10'h223 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h223] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h223]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h223]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h223] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h223]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h224] = (10'h224 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h224] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h224]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h224]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h224] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h224]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h225] = (10'h225 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h225] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h225]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h225]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h225] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h225]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h226] = (10'h226 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h226] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h226]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h226]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h226] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h226]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h227] = (10'h227 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h227] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h227]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h227]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h227] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h227]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h228] = (10'h228 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h228] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h228]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h228]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h228] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h228]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h229] = (10'h229 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h229] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h229]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h229]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h229] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h229]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22a] = (10'h22a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22b] = (10'h22b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22c] = (10'h22c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22d] = (10'h22d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22e] = (10'h22e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22f] = (10'h22f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h230] = (10'h230 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h230] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h230]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h230]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h230] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h230]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h231] = (10'h231 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h231] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h231]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h231]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h231] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h231]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h232] = (10'h232 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h232] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h232]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h232]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h232] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h232]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h233] = (10'h233 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h233] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h233]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h233]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h233] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h233]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h234] = (10'h234 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h234] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h234]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h234]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h234] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h234]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h235] = (10'h235 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h235] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h235]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h235]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h235] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h235]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h236] = (10'h236 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h236] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h236]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h236]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h236] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h236]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h237] = (10'h237 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h237] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h237]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h237]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h237] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h237]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h238] = (10'h238 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h238] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h238]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h238]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h238] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h238]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h239] = (10'h239 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h239] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h239]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h239]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h239] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h239]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23a] = (10'h23a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23b] = (10'h23b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23c] = (10'h23c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23d] = (10'h23d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23e] = (10'h23e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23f] = (10'h23f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h240] = (10'h240 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h240] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h240]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h240]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h240] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h240]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h241] = (10'h241 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h241] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h241]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h241]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h241] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h241]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h242] = (10'h242 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h242] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h242]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h242]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h242] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h242]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h243] = (10'h243 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h243] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h243]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h243]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h243] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h243]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h244] = (10'h244 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h244] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h244]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h244]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h244] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h244]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h245] = (10'h245 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h245] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h245]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h245]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h245] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h245]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h246] = (10'h246 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h246] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h246]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h246]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h246] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h246]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h247] = (10'h247 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h247] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h247]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h247]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h247] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h247]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h248] = (10'h248 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h248] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h248]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h248]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h248] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h248]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h249] = (10'h249 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h249] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h249]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h249]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h249] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h249]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24a] = (10'h24a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24b] = (10'h24b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24c] = (10'h24c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24d] = (10'h24d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24e] = (10'h24e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24f] = (10'h24f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h250] = (10'h250 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h250] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h250]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h250]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h250] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h250]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h251] = (10'h251 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h251] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h251]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h251]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h251] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h251]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h252] = (10'h252 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h252] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h252]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h252]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h252] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h252]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h253] = (10'h253 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h253] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h253]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h253]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h253] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h253]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h254] = (10'h254 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h254] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h254]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h254]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h254] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h254]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h255] = (10'h255 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h255] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h255]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h255]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h255] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h255]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h256] = (10'h256 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h256] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h256]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h256]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h256] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h256]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h257] = (10'h257 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h257] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h257]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h257]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h257] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h257]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h258] = (10'h258 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h258] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h258]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h258]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h258] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h258]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h259] = (10'h259 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h259] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h259]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h259]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h259] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h259]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25a] = (10'h25a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25b] = (10'h25b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25c] = (10'h25c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25d] = (10'h25d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25e] = (10'h25e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25f] = (10'h25f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h260] = (10'h260 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h260] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h260]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h260]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h260] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h260]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h261] = (10'h261 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h261] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h261]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h261]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h261] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h261]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h262] = (10'h262 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h262] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h262]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h262]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h262] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h262]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h263] = (10'h263 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h263] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h263]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h263]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h263] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h263]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h264] = (10'h264 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h264] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h264]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h264]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h264] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h264]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h265] = (10'h265 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h265] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h265]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h265]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h265] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h265]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h266] = (10'h266 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h266] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h266]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h266]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h266] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h266]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h267] = (10'h267 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h267] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h267]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h267]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h267] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h267]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h268] = (10'h268 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h268] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h268]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h268]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h268] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h268]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h269] = (10'h269 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h269] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h269]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h269]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h269] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h269]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26a] = (10'h26a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26b] = (10'h26b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26c] = (10'h26c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26d] = (10'h26d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26e] = (10'h26e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26f] = (10'h26f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h270] = (10'h270 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h270] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h270]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h270]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h270] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h270]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h271] = (10'h271 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h271] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h271]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h271]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h271] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h271]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h272] = (10'h272 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h272] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h272]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h272]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h272] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h272]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h273] = (10'h273 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h273] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h273]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h273]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h273] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h273]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h274] = (10'h274 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h274] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h274]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h274]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h274] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h274]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h275] = (10'h275 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h275] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h275]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h275]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h275] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h275]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h276] = (10'h276 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h276] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h276]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h276]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h276] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h276]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h277] = (10'h277 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h277] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h277]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h277]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h277] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h277]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h278] = (10'h278 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h278] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h278]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h278]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h278] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h278]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h279] = (10'h279 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h279] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h279]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h279]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h279] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h279]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27a] = (10'h27a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27b] = (10'h27b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27c] = (10'h27c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27d] = (10'h27d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27e] = (10'h27e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27f] = (10'h27f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h280] = (10'h280 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h280] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h280]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h280]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h280] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h280]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h281] = (10'h281 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h281] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h281]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h281]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h281] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h281]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h282] = (10'h282 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h282] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h282]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h282]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h282] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h282]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h283] = (10'h283 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h283] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h283]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h283]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h283] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h283]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h284] = (10'h284 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h284] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h284]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h284]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h284] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h284]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h285] = (10'h285 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h285] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h285]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h285]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h285] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h285]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h286] = (10'h286 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h286] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h286]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h286]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h286] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h286]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h287] = (10'h287 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h287] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h287]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h287]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h287] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h287]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h288] = (10'h288 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h288] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h288]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h288]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h288] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h288]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h289] = (10'h289 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h289] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h289]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h289]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h289] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h289]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28a] = (10'h28a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28b] = (10'h28b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28c] = (10'h28c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28d] = (10'h28d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28e] = (10'h28e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28f] = (10'h28f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h290] = (10'h290 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h290] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h290]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h290]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h290] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h290]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h291] = (10'h291 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h291] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h291]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h291]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h291] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h291]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h292] = (10'h292 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h292] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h292]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h292]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h292] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h292]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h293] = (10'h293 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h293] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h293]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h293]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h293] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h293]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h294] = (10'h294 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h294] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h294]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h294]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h294] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h294]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h295] = (10'h295 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h295] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h295]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h295]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h295] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h295]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h296] = (10'h296 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h296] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h296]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h296]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h296] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h296]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h297] = (10'h297 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h297] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h297]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h297]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h297] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h297]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h298] = (10'h298 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h298] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h298]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h298]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h298] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h298]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h299] = (10'h299 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h299] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h299]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h299]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h299] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h299]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29a] = (10'h29a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29b] = (10'h29b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29c] = (10'h29c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29d] = (10'h29d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29e] = (10'h29e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29f] = (10'h29f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a0] = (10'h2a0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a1] = (10'h2a1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a2] = (10'h2a2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a3] = (10'h2a3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a4] = (10'h2a4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a5] = (10'h2a5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a6] = (10'h2a6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a7] = (10'h2a7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a8] = (10'h2a8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a9] = (10'h2a9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2aa] = (10'h2aa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2aa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2aa]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2aa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2aa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2aa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ab] = (10'h2ab == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ab] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ab]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ab]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ab] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ab]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ac] = (10'h2ac == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ac] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ac]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ac]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ac] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ac]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ad] = (10'h2ad == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ad] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ad]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ad]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ad] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ad]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ae] = (10'h2ae == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ae] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ae]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ae]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ae] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ae]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2af] = (10'h2af == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2af] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2af]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2af]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2af] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2af]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b0] = (10'h2b0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b1] = (10'h2b1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b2] = (10'h2b2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b3] = (10'h2b3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b4] = (10'h2b4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b5] = (10'h2b5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b6] = (10'h2b6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b7] = (10'h2b7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b8] = (10'h2b8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b9] = (10'h2b9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ba] = (10'h2ba == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ba] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ba]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ba]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ba] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ba]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bb] = (10'h2bb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bc] = (10'h2bc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bd] = (10'h2bd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2be] = (10'h2be == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2be] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2be]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2be]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2be] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2be]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bf] = (10'h2bf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bf]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c0] = (10'h2c0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c1] = (10'h2c1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c2] = (10'h2c2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c3] = (10'h2c3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c4] = (10'h2c4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c5] = (10'h2c5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c6] = (10'h2c6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c7] = (10'h2c7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c8] = (10'h2c8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c9] = (10'h2c9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ca] = (10'h2ca == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ca] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ca]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ca]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ca] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ca]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cb] = (10'h2cb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cc] = (10'h2cc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cd] = (10'h2cd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ce] = (10'h2ce == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ce] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ce]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ce]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ce] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ce]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cf] = (10'h2cf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cf]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d0] = (10'h2d0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d1] = (10'h2d1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d2] = (10'h2d2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d3] = (10'h2d3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d4] = (10'h2d4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d5] = (10'h2d5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d6] = (10'h2d6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d7] = (10'h2d7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d8] = (10'h2d8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d9] = (10'h2d9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2da] = (10'h2da == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2da] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2da]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2da]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2da] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2da]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2db] = (10'h2db == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2db] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2db]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2db]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2db] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2db]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2dc] = (10'h2dc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2dc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2dc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2dc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2dc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2dc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2dd] = (10'h2dd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2dd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2dd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2dd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2dd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2dd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2de] = (10'h2de == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2de] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2de]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2de]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2de] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2de]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2df] = (10'h2df == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2df] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2df]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2df]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2df] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2df]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e0] = (10'h2e0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e1] = (10'h2e1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e2] = (10'h2e2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e3] = (10'h2e3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e4] = (10'h2e4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e5] = (10'h2e5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e6] = (10'h2e6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e7] = (10'h2e7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e8] = (10'h2e8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e9] = (10'h2e9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ea] = (10'h2ea == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ea] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ea]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ea]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ea] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ea]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2eb] = (10'h2eb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2eb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2eb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2eb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2eb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2eb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ec] = (10'h2ec == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ec] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ec]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ec]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ec] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ec]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ed] = (10'h2ed == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ed] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ed]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ed]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ed] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ed]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ee] = (10'h2ee == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ee] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ee]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ee]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ee] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ee]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ef] = (10'h2ef == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ef] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ef]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ef]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ef] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ef]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f0] = (10'h2f0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f1] = (10'h2f1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f2] = (10'h2f2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f3] = (10'h2f3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f4] = (10'h2f4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f5] = (10'h2f5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f6] = (10'h2f6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f7] = (10'h2f7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f8] = (10'h2f8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f9] = (10'h2f9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fa] = (10'h2fa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fa]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fb] = (10'h2fb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fc] = (10'h2fc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fd] = (10'h2fd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fe] = (10'h2fe == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fe] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fe]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fe]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fe] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fe]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ff] = (10'h2ff == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ff] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ff]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ff]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ff] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ff]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h300] = (10'h300 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h300] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h300]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h300]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h300] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h300]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h301] = (10'h301 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h301] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h301]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h301]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h301] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h301]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h302] = (10'h302 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h302] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h302]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h302]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h302] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h302]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h303] = (10'h303 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h303] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h303]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h303]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h303] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h303]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h304] = (10'h304 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h304] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h304]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h304]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h304] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h304]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h305] = (10'h305 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h305] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h305]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h305]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h305] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h305]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h306] = (10'h306 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h306] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h306]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h306]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h306] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h306]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h307] = (10'h307 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h307] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h307]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h307]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h307] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h307]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h308] = (10'h308 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h308] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h308]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h308]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h308] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h308]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h309] = (10'h309 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h309] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h309]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h309]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h309] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h309]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30a] = (10'h30a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30b] = (10'h30b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30c] = (10'h30c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30d] = (10'h30d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30e] = (10'h30e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30f] = (10'h30f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h310] = (10'h310 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h310] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h310]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h310]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h310] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h310]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h311] = (10'h311 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h311] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h311]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h311]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h311] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h311]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h312] = (10'h312 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h312] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h312]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h312]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h312] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h312]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h313] = (10'h313 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h313] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h313]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h313]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h313] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h313]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h314] = (10'h314 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h314] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h314]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h314]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h314] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h314]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h315] = (10'h315 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h315] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h315]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h315]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h315] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h315]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h316] = (10'h316 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h316] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h316]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h316]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h316] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h316]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h317] = (10'h317 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h317] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h317]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h317]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h317] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h317]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h318] = (10'h318 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h318] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h318]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h318]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h318] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h318]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h319] = (10'h319 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h319] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h319]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h319]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h319] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h319]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31a] = (10'h31a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31b] = (10'h31b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31c] = (10'h31c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31d] = (10'h31d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31e] = (10'h31e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31f] = (10'h31f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h320] = (10'h320 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h320] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h320]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h320]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h320] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h320]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h321] = (10'h321 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h321] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h321]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h321]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h321] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h321]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h322] = (10'h322 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h322] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h322]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h322]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h322] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h322]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h323] = (10'h323 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h323] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h323]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h323]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h323] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h323]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h324] = (10'h324 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h324] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h324]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h324]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h324] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h324]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h325] = (10'h325 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h325] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h325]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h325]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h325] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h325]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h326] = (10'h326 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h326] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h326]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h326]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h326] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h326]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h327] = (10'h327 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h327] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h327]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h327]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h327] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h327]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h328] = (10'h328 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h328] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h328]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h328]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h328] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h328]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h329] = (10'h329 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h329] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h329]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h329]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h329] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h329]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32a] = (10'h32a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32b] = (10'h32b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32c] = (10'h32c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32d] = (10'h32d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32e] = (10'h32e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32f] = (10'h32f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h330] = (10'h330 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h330] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h330]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h330]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h330] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h330]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h331] = (10'h331 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h331] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h331]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h331]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h331] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h331]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h332] = (10'h332 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h332] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h332]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h332]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h332] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h332]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h333] = (10'h333 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h333] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h333]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h333]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h333] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h333]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h334] = (10'h334 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h334] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h334]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h334]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h334] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h334]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h335] = (10'h335 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h335] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h335]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h335]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h335] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h335]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h336] = (10'h336 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h336] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h336]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h336]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h336] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h336]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h337] = (10'h337 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h337] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h337]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h337]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h337] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h337]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h338] = (10'h338 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h338] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h338]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h338]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h338] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h338]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h339] = (10'h339 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h339] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h339]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h339]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h339] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h339]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33a] = (10'h33a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33b] = (10'h33b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33c] = (10'h33c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33d] = (10'h33d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33e] = (10'h33e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33f] = (10'h33f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h340] = (10'h340 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h340] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h340]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h340]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h340] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h340]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h341] = (10'h341 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h341] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h341]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h341]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h341] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h341]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h342] = (10'h342 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h342] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h342]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h342]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h342] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h342]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h343] = (10'h343 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h343] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h343]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h343]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h343] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h343]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h344] = (10'h344 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h344] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h344]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h344]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h344] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h344]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h345] = (10'h345 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h345] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h345]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h345]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h345] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h345]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h346] = (10'h346 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h346] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h346]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h346]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h346] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h346]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h347] = (10'h347 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h347] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h347]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h347]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h347] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h347]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h348] = (10'h348 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h348] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h348]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h348]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h348] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h348]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h349] = (10'h349 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h349] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h349]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h349]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h349] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h349]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34a] = (10'h34a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34b] = (10'h34b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34c] = (10'h34c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34d] = (10'h34d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34e] = (10'h34e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34f] = (10'h34f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h350] = (10'h350 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h350] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h350]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h350]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h350] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h350]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h351] = (10'h351 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h351] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h351]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h351]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h351] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h351]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h352] = (10'h352 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h352] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h352]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h352]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h352] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h352]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h353] = (10'h353 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h353] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h353]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h353]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h353] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h353]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h354] = (10'h354 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h354] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h354]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h354]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h354] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h354]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h355] = (10'h355 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h355] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h355]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h355]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h355] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h355]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h356] = (10'h356 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h356] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h356]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h356]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h356] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h356]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h357] = (10'h357 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h357] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h357]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h357]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h357] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h357]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h358] = (10'h358 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h358] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h358]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h358]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h358] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h358]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h359] = (10'h359 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h359] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h359]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h359]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h359] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h359]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35a] = (10'h35a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35b] = (10'h35b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35c] = (10'h35c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35d] = (10'h35d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35e] = (10'h35e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35f] = (10'h35f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h360] = (10'h360 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h360] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h360]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h360]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h360] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h360]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h361] = (10'h361 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h361] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h361]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h361]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h361] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h361]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h362] = (10'h362 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h362] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h362]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h362]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h362] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h362]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h363] = (10'h363 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h363] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h363]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h363]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h363] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h363]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h364] = (10'h364 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h364] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h364]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h364]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h364] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h364]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h365] = (10'h365 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h365] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h365]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h365]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h365] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h365]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h366] = (10'h366 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h366] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h366]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h366]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h366] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h366]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h367] = (10'h367 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h367] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h367]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h367]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h367] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h367]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h368] = (10'h368 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h368] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h368]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h368]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h368] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h368]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h369] = (10'h369 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h369] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h369]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h369]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h369] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h369]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36a] = (10'h36a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36b] = (10'h36b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36c] = (10'h36c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36d] = (10'h36d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36e] = (10'h36e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36f] = (10'h36f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h370] = (10'h370 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h370] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h370]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h370]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h370] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h370]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h371] = (10'h371 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h371] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h371]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h371]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h371] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h371]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h372] = (10'h372 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h372] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h372]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h372]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h372] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h372]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h373] = (10'h373 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h373] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h373]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h373]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h373] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h373]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h374] = (10'h374 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h374] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h374]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h374]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h374] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h374]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h375] = (10'h375 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h375] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h375]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h375]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h375] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h375]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h376] = (10'h376 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h376] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h376]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h376]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h376] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h376]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h377] = (10'h377 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h377] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h377]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h377]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h377] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h377]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h378] = (10'h378 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h378] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h378]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h378]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h378] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h378]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h379] = (10'h379 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h379] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h379]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h379]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h379] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h379]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37a] = (10'h37a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37b] = (10'h37b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37c] = (10'h37c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37d] = (10'h37d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37e] = (10'h37e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37f] = (10'h37f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h380] = (10'h380 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h380] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h380]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h380]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h380] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h380]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h381] = (10'h381 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h381] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h381]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h381]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h381] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h381]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h382] = (10'h382 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h382] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h382]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h382]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h382] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h382]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h383] = (10'h383 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h383] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h383]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h383]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h383] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h383]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h384] = (10'h384 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h384] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h384]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h384]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h384] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h384]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h385] = (10'h385 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h385] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h385]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h385]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h385] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h385]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h386] = (10'h386 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h386] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h386]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h386]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h386] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h386]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h387] = (10'h387 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h387] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h387]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h387]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h387] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h387]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h388] = (10'h388 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h388] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h388]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h388]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h388] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h388]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h389] = (10'h389 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h389] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h389]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h389]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h389] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h389]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38a] = (10'h38a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38b] = (10'h38b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38c] = (10'h38c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38d] = (10'h38d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38e] = (10'h38e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38f] = (10'h38f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h390] = (10'h390 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h390] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h390]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h390]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h390] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h390]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h391] = (10'h391 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h391] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h391]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h391]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h391] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h391]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h392] = (10'h392 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h392] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h392]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h392]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h392] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h392]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h393] = (10'h393 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h393] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h393]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h393]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h393] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h393]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h394] = (10'h394 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h394] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h394]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h394]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h394] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h394]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h395] = (10'h395 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h395] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h395]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h395]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h395] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h395]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h396] = (10'h396 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h396] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h396]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h396]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h396] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h396]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h397] = (10'h397 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h397] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h397]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h397]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h397] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h397]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h398] = (10'h398 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h398] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h398]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h398]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h398] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h398]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h399] = (10'h399 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h399] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h399]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h399]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h399] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h399]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39a] = (10'h39a == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39a] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39a]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39a]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39a] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39a]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39b] = (10'h39b == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39b] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39b]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39b]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39b] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39b]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39c] = (10'h39c == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39c] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39c]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39c]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39c] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39c]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39d] = (10'h39d == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39d] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39d]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39d]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39d] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39d]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39e] = (10'h39e == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39e] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39e]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39e]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39e] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39e]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39f] = (10'h39f == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39f] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39f]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39f]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39f] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39f]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a0] = (10'h3a0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a1] = (10'h3a1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a2] = (10'h3a2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a3] = (10'h3a3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a4] = (10'h3a4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a5] = (10'h3a5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a6] = (10'h3a6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a7] = (10'h3a7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a8] = (10'h3a8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a9] = (10'h3a9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3aa] = (10'h3aa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3aa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3aa]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3aa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3aa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3aa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ab] = (10'h3ab == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ab] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ab]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ab]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ab] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ab]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ac] = (10'h3ac == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ac] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ac]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ac]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ac] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ac]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ad] = (10'h3ad == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ad] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ad]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ad]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ad] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ad]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ae] = (10'h3ae == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ae] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ae]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ae]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ae] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ae]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3af] = (10'h3af == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3af] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3af]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3af]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3af] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3af]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b0] = (10'h3b0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b1] = (10'h3b1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b2] = (10'h3b2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b3] = (10'h3b3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b4] = (10'h3b4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b5] = (10'h3b5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b6] = (10'h3b6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b7] = (10'h3b7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b8] = (10'h3b8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b9] = (10'h3b9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ba] = (10'h3ba == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ba] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ba]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ba]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ba] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ba]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bb] = (10'h3bb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bc] = (10'h3bc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bd] = (10'h3bd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3be] = (10'h3be == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3be] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3be]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3be]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3be] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3be]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bf] = (10'h3bf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bf]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c0] = (10'h3c0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c1] = (10'h3c1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c2] = (10'h3c2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c3] = (10'h3c3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c4] = (10'h3c4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c5] = (10'h3c5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c6] = (10'h3c6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c7] = (10'h3c7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c8] = (10'h3c8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c9] = (10'h3c9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ca] = (10'h3ca == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ca] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ca]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ca]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ca] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ca]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cb] = (10'h3cb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cc] = (10'h3cc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cd] = (10'h3cd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ce] = (10'h3ce == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ce] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ce]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ce]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ce] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ce]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cf] = (10'h3cf == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cf] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cf]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cf]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cf] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cf]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d0] = (10'h3d0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d1] = (10'h3d1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d2] = (10'h3d2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d3] = (10'h3d3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d4] = (10'h3d4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d5] = (10'h3d5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d6] = (10'h3d6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d7] = (10'h3d7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d8] = (10'h3d8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d9] = (10'h3d9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3da] = (10'h3da == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3da] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3da]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3da]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3da] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3da]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3db] = (10'h3db == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3db] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3db]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3db]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3db] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3db]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3dc] = (10'h3dc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3dc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3dc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3dc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3dc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3dc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3dd] = (10'h3dd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3dd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3dd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3dd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3dd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3dd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3de] = (10'h3de == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3de] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3de]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3de]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3de] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3de]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3df] = (10'h3df == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3df] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3df]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3df]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3df] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3df]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e0] = (10'h3e0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e1] = (10'h3e1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e2] = (10'h3e2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e3] = (10'h3e3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e4] = (10'h3e4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e5] = (10'h3e5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e6] = (10'h3e6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e7] = (10'h3e7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e8] = (10'h3e8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e9] = (10'h3e9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ea] = (10'h3ea == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ea] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ea]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ea]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ea] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ea]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3eb] = (10'h3eb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3eb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3eb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3eb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3eb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3eb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ec] = (10'h3ec == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ec] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ec]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ec]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ec] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ec]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ed] = (10'h3ed == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ed] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ed]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ed]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ed] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ed]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ee] = (10'h3ee == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ee] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ee]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ee]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ee] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ee]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ef] = (10'h3ef == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ef] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ef]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ef]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ef] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ef]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f0] = (10'h3f0 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f0] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f0]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f0]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f0]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f1] = (10'h3f1 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f1] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f1]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f1]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f1] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f1]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f2] = (10'h3f2 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f2] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f2]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f2]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f2] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f2]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f3] = (10'h3f3 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f3] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f3]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f3]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f3] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f3]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f4] = (10'h3f4 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f4] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f4]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f4]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f4] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f4]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f5] = (10'h3f5 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f5] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f5]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f5]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f5] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f5]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f6] = (10'h3f6 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f6] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f6]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f6]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f6] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f6]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f7] = (10'h3f7 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f7] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f7]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f7]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f7] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f7]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f8] = (10'h3f8 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f8] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f8]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f8]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f8] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f8]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f9] = (10'h3f9 == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f9] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f9]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f9]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f9] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f9]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fa] = (10'h3fa == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fa] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fa]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fa]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fa] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fa]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fb] = (10'h3fb == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fb] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fb]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fb]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fb] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fb]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fc] = (10'h3fc == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fc] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fc]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fc]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fc] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fc]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fd] = (10'h3fd == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fd] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fd]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fd]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fd] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fd]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fe] = (10'h3fe == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fe] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fe]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fe]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fe] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fe]));
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ff] = (10'h3ff == axis_fifo_inst__DOT__rd_addr_reg[9:0]) & axis_fifo_inst__DOT__read;
  assign axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ff] = (rst | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ff]) ? (1'b1) : (
                                                                           (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ff]) ? (1'b0) : (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ff] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ff]));
  assign s_axis_tdata__VALID__ = s_axis_tvalid;

  always @(posedge clk) begin
    axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV_Q__ <= axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AV__;
    axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AI_Q__ <= axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____AI__;
    axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____ASSIGN_Q__ <= axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____ASSIGN__;
    axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____VALID_Q__ <= axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____VALID__;
    axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV_Q__ <= axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AV__;
    axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AI_Q__ <= axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____AI__;
    axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN_Q__ <= axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN__;
    axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____VALID_Q__ <= axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____VALID__;
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h40] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h40];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h40] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h40];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h40] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h40];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h40] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h40];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h41] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h41];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h41] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h41];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h41] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h41];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h41] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h41];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h42] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h42];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h42] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h42];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h42] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h42];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h42] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h42];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h43] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h43];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h43] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h43];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h43] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h43];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h43] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h43];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h44] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h44];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h44] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h44];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h44] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h44];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h44] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h44];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h45] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h45];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h45] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h45];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h45] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h45];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h45] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h45];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h46] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h46];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h46] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h46];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h46] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h46];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h46] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h46];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h47] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h47];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h47] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h47];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h47] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h47];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h47] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h47];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h48] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h48];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h48] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h48];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h48] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h48];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h48] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h48];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h49] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h49];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h49] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h49];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h49] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h49];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h49] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h49];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h4f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h4f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h4f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h4f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h4f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h4f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h4f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h4f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h50] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h50];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h50] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h50];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h50] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h50];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h50] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h50];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h51] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h51];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h51] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h51];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h51] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h51];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h51] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h51];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h52] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h52];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h52] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h52];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h52] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h52];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h52] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h52];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h53] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h53];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h53] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h53];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h53] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h53];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h53] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h53];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h54] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h54];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h54] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h54];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h54] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h54];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h54] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h54];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h55] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h55];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h55] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h55];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h55] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h55];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h55] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h55];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h56] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h56];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h56] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h56];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h56] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h56];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h56] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h56];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h57] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h57];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h57] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h57];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h57] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h57];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h57] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h57];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h58] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h58];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h58] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h58];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h58] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h58];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h58] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h58];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h59] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h59];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h59] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h59];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h59] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h59];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h59] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h59];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h5f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h5f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h5f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h5f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h5f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h5f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h5f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h5f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h60] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h60];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h60] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h60];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h60] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h60];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h60] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h60];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h61] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h61];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h61] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h61];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h61] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h61];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h61] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h61];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h62] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h62];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h62] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h62];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h62] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h62];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h62] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h62];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h63] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h63];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h63] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h63];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h63] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h63];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h63] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h63];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h64] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h64];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h64] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h64];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h64] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h64];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h64] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h64];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h65] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h65];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h65] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h65];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h65] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h65];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h65] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h65];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h66] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h66];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h66] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h66];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h66] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h66];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h66] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h66];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h67] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h67];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h67] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h67];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h67] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h67];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h67] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h67];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h68] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h68];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h68] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h68];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h68] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h68];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h68] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h68];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h69] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h69];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h69] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h69];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h69] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h69];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h69] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h69];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h6f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h6f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h6f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h6f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h6f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h6f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h6f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h6f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h70] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h70];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h70] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h70];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h70] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h70];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h70] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h70];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h71] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h71];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h71] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h71];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h71] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h71];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h71] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h71];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h72] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h72];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h72] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h72];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h72] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h72];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h72] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h72];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h73] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h73];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h73] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h73];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h73] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h73];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h73] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h73];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h74] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h74];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h74] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h74];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h74] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h74];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h74] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h74];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h75] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h75];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h75] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h75];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h75] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h75];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h75] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h75];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h76] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h76];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h76] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h76];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h76] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h76];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h76] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h76];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h77] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h77];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h77] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h77];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h77] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h77];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h77] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h77];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h78] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h78];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h78] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h78];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h78] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h78];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h78] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h78];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h79] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h79];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h79] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h79];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h79] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h79];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h79] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h79];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h7f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h7f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h7f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h7f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h7f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h7f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h7f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h7f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h80] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h80];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h80] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h80];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h80] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h80];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h80] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h80];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h81] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h81];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h81] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h81];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h81] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h81];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h81] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h81];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h82] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h82];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h82] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h82];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h82] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h82];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h82] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h82];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h83] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h83];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h83] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h83];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h83] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h83];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h83] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h83];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h84] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h84];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h84] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h84];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h84] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h84];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h84] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h84];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h85] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h85];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h85] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h85];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h85] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h85];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h85] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h85];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h86] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h86];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h86] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h86];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h86] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h86];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h86] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h86];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h87] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h87];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h87] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h87];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h87] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h87];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h87] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h87];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h88] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h88];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h88] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h88];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h88] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h88];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h88] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h88];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h89] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h89];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h89] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h89];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h89] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h89];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h89] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h89];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h8f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h8f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h8f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h8f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h8f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h8f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h8f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h8f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h90] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h90];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h90] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h90];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h90] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h90];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h90] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h90];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h91] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h91];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h91] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h91];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h91] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h91];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h91] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h91];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h92] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h92];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h92] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h92];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h92] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h92];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h92] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h92];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h93] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h93];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h93] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h93];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h93] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h93];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h93] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h93];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h94] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h94];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h94] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h94];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h94] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h94];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h94] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h94];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h95] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h95];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h95] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h95];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h95] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h95];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h95] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h95];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h96] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h96];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h96] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h96];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h96] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h96];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h96] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h96];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h97] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h97];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h97] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h97];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h97] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h97];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h97] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h97];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h98] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h98];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h98] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h98];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h98] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h98];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h98] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h98];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h99] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h99];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h99] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h99];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h99] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h99];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h99] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h99];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h9f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h9f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h9f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h9f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h9f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h9f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h9f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h9f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'ha9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'ha9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'ha9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'ha9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'ha9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'ha9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'ha9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'ha9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'haa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'haa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'haa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'haa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'haa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'haa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'haa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'haa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'had] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'had];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'had] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'had];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'had] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'had];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'had] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'had];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'haf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'haf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'haf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'haf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'haf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'haf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'haf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'haf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hb9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hb9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hb9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hb9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hb9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hb9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hb9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hb9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hbf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hbf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hbf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hbf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hbf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hbf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hbf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hbf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hc9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hc9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hc9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hc9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hc9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hc9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hc9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hc9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hcf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hcf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hcf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hcf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hcf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hcf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hcf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hcf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hd9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hd9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hd9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hd9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hd9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hd9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hd9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hd9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hda] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hda];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hda] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hda];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hda] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hda];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hda] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hda];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hde] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hde];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hde] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hde];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hde] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hde];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hde] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hde];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hdf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hdf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hdf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hdf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hdf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hdf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hdf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hdf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'he9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'he9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'he9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'he9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'he9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'he9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'he9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'he9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'heb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'heb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'heb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'heb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'heb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'heb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'heb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'heb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hf9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hf9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hf9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hf9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hf9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hf9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hf9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hf9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hfe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hfe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hfe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hfe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hfe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hfe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hfe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hfe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'hff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'hff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'hff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'hff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'hff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'hff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'hff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'hff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h100] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h100];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h100] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h100];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h100] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h100];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h100] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h100];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h101] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h101];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h101] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h101];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h101] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h101];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h101] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h101];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h102] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h102];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h102] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h102];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h102] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h102];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h102] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h102];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h103] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h103];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h103] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h103];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h103] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h103];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h103] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h103];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h104] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h104];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h104] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h104];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h104] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h104];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h104] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h104];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h105] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h105];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h105] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h105];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h105] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h105];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h105] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h105];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h106] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h106];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h106] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h106];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h106] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h106];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h106] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h106];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h107] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h107];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h107] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h107];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h107] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h107];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h107] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h107];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h108] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h108];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h108] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h108];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h108] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h108];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h108] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h108];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h109] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h109];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h109] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h109];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h109] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h109];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h109] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h109];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h10f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h10f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h10f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h10f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h10f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h10f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h10f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h10f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h110] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h110];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h110] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h110];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h110] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h110];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h110] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h110];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h111] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h111];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h111] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h111];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h111] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h111];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h111] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h111];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h112] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h112];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h112] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h112];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h112] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h112];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h112] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h112];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h113] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h113];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h113] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h113];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h113] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h113];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h113] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h113];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h114] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h114];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h114] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h114];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h114] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h114];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h114] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h114];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h115] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h115];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h115] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h115];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h115] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h115];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h115] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h115];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h116] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h116];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h116] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h116];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h116] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h116];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h116] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h116];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h117] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h117];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h117] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h117];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h117] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h117];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h117] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h117];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h118] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h118];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h118] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h118];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h118] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h118];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h118] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h118];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h119] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h119];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h119] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h119];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h119] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h119];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h119] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h119];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h11f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h11f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h11f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h11f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h11f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h11f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h11f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h11f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h120] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h120];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h120] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h120];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h120] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h120];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h120] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h120];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h121] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h121];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h121] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h121];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h121] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h121];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h121] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h121];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h122] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h122];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h122] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h122];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h122] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h122];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h122] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h122];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h123] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h123];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h123] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h123];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h123] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h123];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h123] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h123];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h124] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h124];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h124] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h124];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h124] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h124];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h124] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h124];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h125] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h125];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h125] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h125];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h125] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h125];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h125] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h125];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h126] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h126];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h126] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h126];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h126] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h126];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h126] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h126];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h127] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h127];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h127] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h127];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h127] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h127];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h127] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h127];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h128] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h128];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h128] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h128];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h128] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h128];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h128] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h128];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h129] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h129];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h129] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h129];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h129] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h129];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h129] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h129];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h12f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h12f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h12f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h12f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h12f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h12f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h12f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h12f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h130] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h130];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h130] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h130];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h130] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h130];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h130] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h130];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h131] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h131];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h131] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h131];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h131] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h131];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h131] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h131];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h132] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h132];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h132] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h132];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h132] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h132];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h132] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h132];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h133] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h133];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h133] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h133];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h133] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h133];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h133] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h133];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h134] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h134];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h134] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h134];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h134] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h134];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h134] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h134];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h135] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h135];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h135] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h135];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h135] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h135];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h135] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h135];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h136] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h136];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h136] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h136];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h136] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h136];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h136] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h136];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h137] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h137];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h137] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h137];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h137] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h137];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h137] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h137];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h138] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h138];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h138] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h138];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h138] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h138];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h138] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h138];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h139] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h139];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h139] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h139];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h139] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h139];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h139] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h139];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h13f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h13f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h13f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h13f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h13f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h13f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h13f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h13f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h140] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h140];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h140] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h140];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h140] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h140];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h140] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h140];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h141] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h141];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h141] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h141];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h141] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h141];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h141] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h141];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h142] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h142];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h142] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h142];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h142] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h142];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h142] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h142];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h143] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h143];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h143] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h143];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h143] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h143];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h143] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h143];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h144] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h144];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h144] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h144];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h144] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h144];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h144] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h144];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h145] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h145];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h145] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h145];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h145] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h145];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h145] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h145];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h146] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h146];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h146] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h146];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h146] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h146];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h146] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h146];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h147] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h147];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h147] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h147];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h147] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h147];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h147] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h147];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h148] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h148];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h148] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h148];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h148] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h148];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h148] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h148];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h149] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h149];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h149] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h149];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h149] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h149];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h149] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h149];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h14f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h14f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h14f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h14f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h14f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h14f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h14f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h14f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h150] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h150];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h150] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h150];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h150] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h150];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h150] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h150];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h151] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h151];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h151] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h151];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h151] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h151];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h151] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h151];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h152] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h152];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h152] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h152];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h152] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h152];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h152] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h152];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h153] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h153];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h153] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h153];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h153] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h153];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h153] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h153];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h154] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h154];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h154] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h154];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h154] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h154];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h154] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h154];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h155] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h155];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h155] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h155];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h155] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h155];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h155] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h155];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h156] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h156];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h156] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h156];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h156] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h156];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h156] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h156];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h157] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h157];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h157] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h157];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h157] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h157];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h157] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h157];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h158] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h158];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h158] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h158];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h158] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h158];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h158] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h158];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h159] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h159];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h159] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h159];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h159] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h159];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h159] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h159];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h15f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h15f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h15f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h15f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h15f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h15f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h15f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h15f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h160] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h160];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h160] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h160];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h160] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h160];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h160] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h160];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h161] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h161];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h161] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h161];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h161] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h161];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h161] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h161];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h162] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h162];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h162] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h162];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h162] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h162];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h162] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h162];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h163] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h163];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h163] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h163];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h163] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h163];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h163] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h163];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h164] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h164];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h164] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h164];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h164] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h164];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h164] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h164];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h165] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h165];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h165] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h165];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h165] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h165];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h165] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h165];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h166] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h166];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h166] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h166];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h166] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h166];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h166] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h166];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h167] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h167];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h167] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h167];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h167] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h167];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h167] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h167];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h168] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h168];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h168] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h168];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h168] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h168];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h168] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h168];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h169] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h169];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h169] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h169];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h169] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h169];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h169] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h169];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h16f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h16f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h16f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h16f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h16f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h16f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h16f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h16f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h170] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h170];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h170] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h170];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h170] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h170];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h170] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h170];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h171] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h171];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h171] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h171];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h171] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h171];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h171] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h171];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h172] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h172];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h172] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h172];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h172] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h172];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h172] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h172];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h173] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h173];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h173] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h173];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h173] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h173];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h173] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h173];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h174] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h174];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h174] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h174];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h174] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h174];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h174] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h174];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h175] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h175];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h175] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h175];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h175] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h175];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h175] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h175];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h176] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h176];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h176] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h176];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h176] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h176];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h176] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h176];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h177] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h177];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h177] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h177];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h177] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h177];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h177] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h177];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h178] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h178];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h178] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h178];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h178] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h178];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h178] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h178];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h179] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h179];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h179] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h179];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h179] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h179];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h179] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h179];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h17f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h17f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h17f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h17f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h17f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h17f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h17f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h17f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h180] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h180];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h180] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h180];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h180] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h180];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h180] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h180];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h181] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h181];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h181] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h181];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h181] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h181];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h181] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h181];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h182] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h182];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h182] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h182];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h182] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h182];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h182] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h182];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h183] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h183];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h183] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h183];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h183] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h183];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h183] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h183];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h184] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h184];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h184] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h184];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h184] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h184];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h184] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h184];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h185] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h185];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h185] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h185];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h185] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h185];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h185] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h185];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h186] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h186];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h186] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h186];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h186] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h186];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h186] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h186];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h187] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h187];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h187] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h187];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h187] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h187];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h187] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h187];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h188] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h188];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h188] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h188];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h188] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h188];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h188] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h188];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h189] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h189];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h189] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h189];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h189] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h189];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h189] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h189];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h18f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h18f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h18f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h18f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h18f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h18f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h18f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h18f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h190] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h190];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h190] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h190];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h190] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h190];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h190] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h190];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h191] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h191];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h191] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h191];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h191] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h191];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h191] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h191];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h192] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h192];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h192] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h192];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h192] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h192];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h192] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h192];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h193] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h193];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h193] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h193];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h193] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h193];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h193] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h193];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h194] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h194];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h194] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h194];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h194] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h194];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h194] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h194];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h195] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h195];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h195] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h195];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h195] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h195];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h195] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h195];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h196] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h196];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h196] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h196];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h196] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h196];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h196] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h196];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h197] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h197];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h197] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h197];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h197] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h197];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h197] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h197];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h198] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h198];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h198] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h198];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h198] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h198];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h198] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h198];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h199] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h199];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h199] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h199];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h199] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h199];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h199] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h199];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h19f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h19f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h19f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h19f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h19f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h19f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h19f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h19f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h1ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h1ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h1ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h1ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h1ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h1ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h1ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h1ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h200] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h200];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h200] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h200];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h200] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h200];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h200] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h200];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h201] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h201];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h201] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h201];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h201] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h201];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h201] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h201];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h202] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h202];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h202] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h202];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h202] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h202];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h202] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h202];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h203] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h203];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h203] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h203];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h203] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h203];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h203] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h203];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h204] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h204];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h204] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h204];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h204] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h204];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h204] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h204];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h205] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h205];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h205] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h205];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h205] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h205];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h205] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h205];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h206] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h206];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h206] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h206];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h206] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h206];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h206] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h206];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h207] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h207];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h207] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h207];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h207] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h207];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h207] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h207];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h208] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h208];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h208] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h208];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h208] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h208];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h208] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h208];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h209] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h209];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h209] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h209];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h209] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h209];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h209] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h209];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h20f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h20f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h20f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h20f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h20f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h20f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h20f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h20f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h210] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h210];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h210] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h210];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h210] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h210];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h210] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h210];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h211] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h211];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h211] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h211];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h211] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h211];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h211] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h211];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h212] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h212];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h212] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h212];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h212] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h212];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h212] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h212];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h213] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h213];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h213] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h213];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h213] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h213];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h213] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h213];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h214] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h214];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h214] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h214];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h214] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h214];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h214] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h214];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h215] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h215];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h215] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h215];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h215] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h215];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h215] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h215];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h216] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h216];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h216] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h216];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h216] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h216];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h216] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h216];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h217] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h217];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h217] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h217];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h217] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h217];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h217] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h217];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h218] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h218];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h218] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h218];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h218] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h218];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h218] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h218];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h219] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h219];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h219] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h219];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h219] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h219];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h219] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h219];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h21f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h21f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h21f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h21f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h21f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h21f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h21f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h21f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h220] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h220];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h220] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h220];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h220] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h220];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h220] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h220];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h221] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h221];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h221] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h221];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h221] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h221];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h221] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h221];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h222] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h222];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h222] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h222];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h222] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h222];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h222] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h222];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h223] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h223];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h223] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h223];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h223] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h223];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h223] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h223];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h224] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h224];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h224] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h224];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h224] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h224];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h224] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h224];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h225] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h225];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h225] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h225];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h225] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h225];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h225] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h225];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h226] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h226];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h226] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h226];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h226] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h226];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h226] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h226];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h227] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h227];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h227] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h227];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h227] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h227];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h227] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h227];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h228] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h228];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h228] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h228];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h228] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h228];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h228] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h228];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h229] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h229];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h229] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h229];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h229] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h229];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h229] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h229];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h22f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h22f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h22f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h22f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h22f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h22f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h22f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h22f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h230] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h230];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h230] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h230];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h230] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h230];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h230] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h230];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h231] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h231];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h231] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h231];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h231] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h231];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h231] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h231];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h232] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h232];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h232] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h232];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h232] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h232];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h232] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h232];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h233] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h233];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h233] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h233];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h233] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h233];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h233] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h233];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h234] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h234];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h234] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h234];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h234] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h234];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h234] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h234];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h235] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h235];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h235] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h235];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h235] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h235];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h235] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h235];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h236] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h236];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h236] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h236];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h236] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h236];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h236] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h236];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h237] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h237];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h237] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h237];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h237] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h237];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h237] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h237];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h238] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h238];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h238] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h238];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h238] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h238];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h238] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h238];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h239] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h239];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h239] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h239];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h239] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h239];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h239] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h239];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h23f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h23f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h23f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h23f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h23f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h23f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h23f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h23f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h240] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h240];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h240] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h240];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h240] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h240];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h240] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h240];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h241] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h241];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h241] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h241];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h241] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h241];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h241] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h241];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h242] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h242];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h242] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h242];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h242] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h242];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h242] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h242];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h243] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h243];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h243] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h243];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h243] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h243];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h243] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h243];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h244] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h244];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h244] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h244];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h244] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h244];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h244] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h244];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h245] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h245];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h245] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h245];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h245] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h245];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h245] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h245];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h246] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h246];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h246] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h246];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h246] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h246];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h246] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h246];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h247] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h247];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h247] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h247];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h247] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h247];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h247] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h247];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h248] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h248];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h248] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h248];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h248] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h248];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h248] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h248];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h249] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h249];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h249] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h249];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h249] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h249];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h249] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h249];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h24f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h24f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h24f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h24f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h24f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h24f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h24f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h24f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h250] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h250];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h250] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h250];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h250] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h250];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h250] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h250];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h251] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h251];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h251] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h251];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h251] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h251];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h251] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h251];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h252] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h252];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h252] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h252];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h252] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h252];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h252] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h252];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h253] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h253];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h253] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h253];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h253] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h253];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h253] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h253];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h254] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h254];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h254] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h254];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h254] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h254];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h254] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h254];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h255] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h255];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h255] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h255];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h255] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h255];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h255] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h255];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h256] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h256];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h256] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h256];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h256] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h256];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h256] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h256];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h257] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h257];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h257] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h257];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h257] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h257];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h257] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h257];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h258] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h258];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h258] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h258];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h258] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h258];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h258] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h258];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h259] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h259];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h259] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h259];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h259] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h259];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h259] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h259];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h25f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h25f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h25f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h25f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h25f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h25f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h25f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h25f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h260] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h260];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h260] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h260];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h260] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h260];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h260] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h260];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h261] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h261];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h261] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h261];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h261] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h261];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h261] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h261];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h262] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h262];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h262] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h262];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h262] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h262];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h262] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h262];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h263] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h263];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h263] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h263];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h263] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h263];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h263] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h263];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h264] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h264];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h264] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h264];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h264] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h264];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h264] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h264];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h265] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h265];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h265] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h265];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h265] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h265];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h265] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h265];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h266] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h266];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h266] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h266];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h266] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h266];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h266] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h266];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h267] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h267];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h267] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h267];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h267] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h267];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h267] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h267];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h268] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h268];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h268] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h268];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h268] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h268];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h268] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h268];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h269] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h269];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h269] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h269];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h269] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h269];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h269] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h269];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h26f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h26f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h26f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h26f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h26f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h26f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h26f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h26f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h270] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h270];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h270] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h270];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h270] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h270];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h270] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h270];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h271] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h271];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h271] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h271];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h271] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h271];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h271] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h271];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h272] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h272];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h272] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h272];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h272] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h272];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h272] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h272];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h273] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h273];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h273] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h273];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h273] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h273];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h273] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h273];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h274] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h274];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h274] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h274];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h274] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h274];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h274] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h274];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h275] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h275];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h275] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h275];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h275] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h275];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h275] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h275];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h276] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h276];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h276] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h276];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h276] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h276];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h276] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h276];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h277] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h277];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h277] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h277];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h277] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h277];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h277] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h277];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h278] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h278];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h278] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h278];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h278] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h278];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h278] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h278];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h279] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h279];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h279] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h279];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h279] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h279];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h279] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h279];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h27f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h27f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h27f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h27f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h27f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h27f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h27f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h27f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h280] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h280];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h280] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h280];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h280] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h280];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h280] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h280];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h281] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h281];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h281] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h281];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h281] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h281];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h281] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h281];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h282] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h282];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h282] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h282];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h282] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h282];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h282] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h282];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h283] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h283];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h283] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h283];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h283] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h283];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h283] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h283];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h284] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h284];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h284] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h284];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h284] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h284];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h284] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h284];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h285] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h285];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h285] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h285];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h285] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h285];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h285] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h285];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h286] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h286];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h286] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h286];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h286] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h286];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h286] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h286];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h287] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h287];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h287] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h287];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h287] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h287];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h287] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h287];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h288] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h288];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h288] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h288];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h288] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h288];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h288] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h288];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h289] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h289];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h289] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h289];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h289] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h289];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h289] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h289];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h28f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h28f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h28f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h28f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h28f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h28f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h28f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h28f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h290] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h290];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h290] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h290];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h290] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h290];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h290] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h290];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h291] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h291];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h291] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h291];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h291] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h291];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h291] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h291];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h292] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h292];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h292] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h292];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h292] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h292];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h292] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h292];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h293] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h293];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h293] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h293];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h293] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h293];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h293] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h293];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h294] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h294];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h294] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h294];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h294] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h294];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h294] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h294];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h295] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h295];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h295] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h295];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h295] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h295];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h295] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h295];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h296] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h296];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h296] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h296];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h296] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h296];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h296] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h296];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h297] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h297];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h297] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h297];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h297] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h297];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h297] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h297];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h298] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h298];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h298] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h298];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h298] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h298];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h298] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h298];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h299] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h299];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h299] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h299];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h299] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h299];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h299] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h299];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h29f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h29f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h29f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h29f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h29f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h29f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h29f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h29f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h2ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h2ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h2ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h2ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h2ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h2ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h2ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h2ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h300] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h300];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h300] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h300];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h300] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h300];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h300] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h300];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h301] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h301];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h301] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h301];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h301] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h301];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h301] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h301];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h302] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h302];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h302] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h302];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h302] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h302];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h302] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h302];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h303] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h303];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h303] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h303];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h303] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h303];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h303] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h303];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h304] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h304];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h304] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h304];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h304] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h304];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h304] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h304];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h305] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h305];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h305] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h305];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h305] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h305];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h305] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h305];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h306] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h306];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h306] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h306];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h306] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h306];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h306] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h306];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h307] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h307];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h307] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h307];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h307] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h307];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h307] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h307];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h308] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h308];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h308] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h308];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h308] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h308];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h308] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h308];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h309] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h309];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h309] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h309];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h309] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h309];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h309] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h309];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h30f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h30f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h30f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h30f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h30f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h30f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h30f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h30f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h310] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h310];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h310] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h310];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h310] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h310];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h310] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h310];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h311] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h311];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h311] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h311];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h311] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h311];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h311] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h311];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h312] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h312];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h312] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h312];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h312] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h312];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h312] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h312];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h313] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h313];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h313] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h313];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h313] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h313];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h313] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h313];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h314] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h314];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h314] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h314];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h314] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h314];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h314] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h314];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h315] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h315];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h315] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h315];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h315] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h315];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h315] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h315];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h316] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h316];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h316] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h316];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h316] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h316];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h316] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h316];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h317] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h317];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h317] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h317];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h317] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h317];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h317] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h317];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h318] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h318];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h318] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h318];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h318] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h318];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h318] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h318];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h319] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h319];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h319] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h319];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h319] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h319];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h319] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h319];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h31f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h31f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h31f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h31f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h31f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h31f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h31f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h31f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h320] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h320];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h320] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h320];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h320] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h320];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h320] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h320];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h321] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h321];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h321] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h321];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h321] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h321];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h321] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h321];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h322] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h322];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h322] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h322];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h322] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h322];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h322] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h322];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h323] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h323];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h323] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h323];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h323] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h323];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h323] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h323];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h324] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h324];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h324] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h324];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h324] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h324];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h324] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h324];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h325] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h325];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h325] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h325];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h325] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h325];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h325] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h325];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h326] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h326];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h326] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h326];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h326] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h326];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h326] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h326];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h327] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h327];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h327] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h327];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h327] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h327];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h327] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h327];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h328] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h328];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h328] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h328];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h328] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h328];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h328] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h328];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h329] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h329];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h329] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h329];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h329] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h329];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h329] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h329];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h32f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h32f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h32f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h32f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h32f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h32f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h32f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h32f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h330] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h330];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h330] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h330];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h330] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h330];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h330] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h330];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h331] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h331];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h331] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h331];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h331] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h331];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h331] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h331];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h332] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h332];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h332] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h332];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h332] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h332];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h332] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h332];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h333] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h333];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h333] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h333];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h333] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h333];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h333] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h333];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h334] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h334];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h334] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h334];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h334] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h334];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h334] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h334];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h335] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h335];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h335] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h335];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h335] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h335];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h335] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h335];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h336] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h336];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h336] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h336];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h336] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h336];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h336] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h336];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h337] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h337];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h337] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h337];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h337] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h337];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h337] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h337];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h338] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h338];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h338] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h338];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h338] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h338];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h338] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h338];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h339] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h339];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h339] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h339];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h339] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h339];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h339] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h339];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h33f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h33f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h33f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h33f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h33f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h33f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h33f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h33f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h340] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h340];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h340] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h340];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h340] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h340];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h340] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h340];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h341] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h341];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h341] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h341];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h341] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h341];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h341] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h341];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h342] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h342];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h342] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h342];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h342] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h342];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h342] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h342];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h343] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h343];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h343] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h343];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h343] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h343];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h343] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h343];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h344] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h344];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h344] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h344];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h344] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h344];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h344] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h344];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h345] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h345];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h345] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h345];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h345] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h345];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h345] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h345];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h346] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h346];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h346] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h346];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h346] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h346];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h346] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h346];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h347] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h347];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h347] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h347];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h347] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h347];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h347] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h347];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h348] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h348];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h348] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h348];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h348] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h348];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h348] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h348];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h349] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h349];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h349] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h349];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h349] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h349];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h349] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h349];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h34f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h34f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h34f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h34f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h34f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h34f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h34f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h34f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h350] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h350];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h350] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h350];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h350] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h350];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h350] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h350];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h351] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h351];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h351] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h351];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h351] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h351];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h351] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h351];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h352] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h352];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h352] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h352];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h352] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h352];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h352] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h352];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h353] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h353];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h353] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h353];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h353] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h353];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h353] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h353];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h354] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h354];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h354] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h354];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h354] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h354];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h354] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h354];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h355] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h355];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h355] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h355];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h355] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h355];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h355] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h355];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h356] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h356];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h356] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h356];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h356] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h356];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h356] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h356];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h357] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h357];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h357] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h357];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h357] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h357];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h357] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h357];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h358] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h358];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h358] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h358];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h358] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h358];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h358] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h358];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h359] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h359];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h359] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h359];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h359] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h359];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h359] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h359];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h35f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h35f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h35f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h35f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h35f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h35f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h35f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h35f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h360] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h360];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h360] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h360];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h360] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h360];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h360] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h360];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h361] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h361];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h361] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h361];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h361] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h361];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h361] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h361];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h362] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h362];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h362] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h362];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h362] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h362];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h362] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h362];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h363] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h363];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h363] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h363];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h363] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h363];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h363] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h363];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h364] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h364];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h364] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h364];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h364] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h364];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h364] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h364];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h365] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h365];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h365] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h365];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h365] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h365];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h365] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h365];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h366] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h366];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h366] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h366];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h366] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h366];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h366] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h366];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h367] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h367];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h367] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h367];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h367] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h367];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h367] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h367];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h368] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h368];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h368] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h368];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h368] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h368];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h368] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h368];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h369] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h369];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h369] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h369];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h369] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h369];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h369] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h369];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h36f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h36f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h36f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h36f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h36f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h36f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h36f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h36f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h370] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h370];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h370] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h370];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h370] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h370];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h370] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h370];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h371] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h371];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h371] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h371];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h371] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h371];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h371] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h371];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h372] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h372];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h372] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h372];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h372] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h372];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h372] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h372];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h373] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h373];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h373] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h373];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h373] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h373];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h373] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h373];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h374] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h374];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h374] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h374];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h374] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h374];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h374] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h374];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h375] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h375];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h375] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h375];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h375] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h375];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h375] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h375];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h376] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h376];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h376] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h376];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h376] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h376];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h376] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h376];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h377] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h377];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h377] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h377];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h377] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h377];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h377] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h377];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h378] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h378];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h378] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h378];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h378] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h378];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h378] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h378];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h379] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h379];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h379] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h379];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h379] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h379];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h379] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h379];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h37f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h37f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h37f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h37f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h37f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h37f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h37f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h37f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h380] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h380];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h380] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h380];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h380] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h380];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h380] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h380];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h381] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h381];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h381] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h381];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h381] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h381];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h381] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h381];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h382] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h382];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h382] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h382];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h382] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h382];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h382] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h382];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h383] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h383];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h383] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h383];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h383] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h383];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h383] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h383];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h384] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h384];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h384] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h384];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h384] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h384];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h384] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h384];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h385] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h385];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h385] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h385];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h385] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h385];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h385] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h385];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h386] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h386];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h386] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h386];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h386] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h386];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h386] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h386];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h387] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h387];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h387] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h387];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h387] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h387];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h387] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h387];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h388] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h388];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h388] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h388];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h388] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h388];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h388] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h388];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h389] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h389];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h389] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h389];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h389] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h389];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h389] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h389];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h38f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h38f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h38f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h38f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h38f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h38f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h38f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h38f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h390] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h390];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h390] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h390];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h390] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h390];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h390] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h390];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h391] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h391];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h391] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h391];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h391] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h391];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h391] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h391];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h392] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h392];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h392] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h392];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h392] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h392];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h392] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h392];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h393] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h393];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h393] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h393];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h393] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h393];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h393] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h393];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h394] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h394];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h394] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h394];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h394] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h394];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h394] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h394];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h395] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h395];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h395] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h395];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h395] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h395];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h395] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h395];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h396] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h396];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h396] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h396];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h396] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h396];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h396] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h396];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h397] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h397];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h397] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h397];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h397] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h397];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h397] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h397];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h398] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h398];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h398] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h398];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h398] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h398];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h398] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h398];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h399] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h399];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h399] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h399];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h399] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h399];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h399] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h399];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h39f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h39f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h39f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h39f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h39f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h39f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h39f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h39f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV_Q__[10'h3ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AV__[10'h3ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI_Q__[10'h3ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____AI__[10'h3ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[10'h3ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN__[10'h3ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID_Q__[10'h3ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____VALID__[10'h3ff];
    axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____PROP_Q__ <= axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____PROP__;
    axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____GOOD_Q__ <= axis_fifo_inst__DOT__m_axis_reg__BRA__31__03A0__KET____GOOD__;
    axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP_Q__ <= axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP__;
    axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD_Q__ <= axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD__;
    if (~(axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD_Q__ | axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP_Q__) & axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN_Q__) $display("[%0t] %%loss: axis_fifo_wrapper.axis_fifo_inst__DOT__mem_read_data_reg 'd31 'd0 None None", $time ) /*debug_display_flowguard*/; 
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h40] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h40];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h40] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h40];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h41] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h41];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h41] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h41];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h42] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h42];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h42] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h42];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h43] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h43];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h43] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h43];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h44] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h44];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h44] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h44];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h45] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h45];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h45] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h45];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h46] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h46];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h46] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h46];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h47] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h47];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h47] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h47];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h48] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h48];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h48] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h48];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h49] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h49];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h49] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h49];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h4f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h4f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h4f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h4f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h50] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h50];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h50] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h50];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h51] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h51];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h51] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h51];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h52] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h52];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h52] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h52];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h53] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h53];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h53] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h53];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h54] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h54];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h54] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h54];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h55] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h55];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h55] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h55];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h56] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h56];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h56] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h56];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h57] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h57];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h57] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h57];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h58] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h58];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h58] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h58];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h59] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h59];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h59] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h59];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h5f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h5f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h5f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h5f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h60] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h60];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h60] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h60];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h61] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h61];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h61] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h61];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h62] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h62];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h62] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h62];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h63] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h63];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h63] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h63];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h64] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h64];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h64] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h64];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h65] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h65];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h65] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h65];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h66] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h66];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h66] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h66];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h67] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h67];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h67] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h67];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h68] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h68];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h68] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h68];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h69] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h69];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h69] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h69];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h6f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h6f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h6f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h6f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h70] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h70];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h70] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h70];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h71] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h71];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h71] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h71];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h72] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h72];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h72] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h72];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h73] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h73];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h73] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h73];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h74] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h74];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h74] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h74];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h75] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h75];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h75] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h75];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h76] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h76];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h76] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h76];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h77] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h77];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h77] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h77];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h78] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h78];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h78] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h78];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h79] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h79];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h79] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h79];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h7f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h7f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h7f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h7f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h80] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h80];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h80] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h80];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h81] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h81];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h81] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h81];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h82] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h82];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h82] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h82];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h83] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h83];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h83] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h83];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h84] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h84];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h84] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h84];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h85] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h85];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h85] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h85];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h86] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h86];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h86] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h86];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h87] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h87];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h87] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h87];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h88] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h88];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h88] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h88];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h89] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h89];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h89] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h89];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h8f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h8f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h8f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h8f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h90] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h90];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h90] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h90];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h91] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h91];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h91] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h91];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h92] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h92];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h92] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h92];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h93] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h93];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h93] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h93];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h94] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h94];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h94] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h94];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h95] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h95];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h95] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h95];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h96] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h96];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h96] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h96];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h97] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h97];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h97] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h97];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h98] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h98];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h98] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h98];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h99] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h99];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h99] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h99];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h9f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h9f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h9f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h9f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'ha9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'ha9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'ha9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'ha9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'haa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'haa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'haa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'haa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'had] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'had];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'had] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'had];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'haf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'haf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'haf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'haf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hb9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hb9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hb9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hb9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hbf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hbf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hbf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hbf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hc9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hc9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hc9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hc9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hcf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hcf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hcf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hcf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hd9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hd9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hd9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hd9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hda] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hda];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hda] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hda];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hde] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hde];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hde] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hde];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hdf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hdf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hdf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hdf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'he9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'he9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'he9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'he9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'heb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'heb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'heb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'heb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hf9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hf9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hf9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hf9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hfe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hfe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hfe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hfe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'hff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'hff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'hff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'hff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h100] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h100];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h100] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h100];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h101] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h101];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h101] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h101];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h102] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h102];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h102] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h102];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h103] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h103];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h103] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h103];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h104] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h104];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h104] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h104];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h105] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h105];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h105] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h105];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h106] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h106];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h106] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h106];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h107] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h107];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h107] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h107];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h108] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h108];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h108] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h108];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h109] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h109];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h109] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h109];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h10f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h10f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h10f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h10f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h110] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h110];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h110] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h110];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h111] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h111];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h111] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h111];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h112] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h112];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h112] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h112];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h113] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h113];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h113] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h113];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h114] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h114];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h114] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h114];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h115] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h115];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h115] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h115];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h116] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h116];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h116] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h116];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h117] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h117];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h117] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h117];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h118] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h118];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h118] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h118];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h119] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h119];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h119] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h119];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h11f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h11f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h11f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h11f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h120] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h120];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h120] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h120];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h121] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h121];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h121] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h121];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h122] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h122];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h122] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h122];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h123] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h123];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h123] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h123];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h124] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h124];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h124] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h124];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h125] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h125];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h125] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h125];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h126] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h126];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h126] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h126];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h127] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h127];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h127] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h127];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h128] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h128];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h128] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h128];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h129] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h129];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h129] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h129];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h12f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h12f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h12f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h12f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h130] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h130];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h130] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h130];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h131] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h131];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h131] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h131];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h132] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h132];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h132] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h132];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h133] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h133];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h133] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h133];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h134] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h134];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h134] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h134];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h135] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h135];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h135] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h135];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h136] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h136];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h136] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h136];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h137] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h137];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h137] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h137];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h138] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h138];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h138] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h138];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h139] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h139];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h139] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h139];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h13f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h13f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h13f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h13f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h140] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h140];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h140] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h140];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h141] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h141];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h141] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h141];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h142] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h142];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h142] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h142];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h143] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h143];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h143] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h143];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h144] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h144];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h144] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h144];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h145] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h145];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h145] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h145];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h146] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h146];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h146] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h146];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h147] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h147];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h147] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h147];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h148] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h148];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h148] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h148];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h149] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h149];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h149] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h149];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h14f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h14f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h14f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h14f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h150] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h150];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h150] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h150];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h151] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h151];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h151] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h151];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h152] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h152];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h152] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h152];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h153] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h153];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h153] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h153];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h154] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h154];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h154] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h154];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h155] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h155];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h155] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h155];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h156] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h156];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h156] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h156];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h157] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h157];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h157] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h157];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h158] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h158];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h158] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h158];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h159] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h159];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h159] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h159];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h15f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h15f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h15f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h15f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h160] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h160];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h160] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h160];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h161] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h161];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h161] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h161];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h162] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h162];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h162] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h162];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h163] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h163];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h163] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h163];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h164] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h164];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h164] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h164];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h165] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h165];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h165] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h165];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h166] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h166];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h166] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h166];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h167] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h167];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h167] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h167];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h168] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h168];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h168] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h168];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h169] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h169];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h169] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h169];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h16f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h16f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h16f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h16f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h170] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h170];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h170] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h170];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h171] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h171];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h171] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h171];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h172] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h172];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h172] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h172];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h173] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h173];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h173] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h173];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h174] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h174];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h174] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h174];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h175] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h175];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h175] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h175];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h176] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h176];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h176] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h176];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h177] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h177];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h177] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h177];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h178] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h178];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h178] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h178];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h179] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h179];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h179] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h179];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h17f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h17f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h17f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h17f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h180] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h180];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h180] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h180];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h181] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h181];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h181] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h181];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h182] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h182];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h182] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h182];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h183] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h183];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h183] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h183];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h184] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h184];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h184] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h184];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h185] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h185];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h185] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h185];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h186] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h186];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h186] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h186];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h187] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h187];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h187] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h187];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h188] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h188];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h188] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h188];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h189] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h189];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h189] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h189];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h18f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h18f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h18f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h18f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h190] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h190];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h190] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h190];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h191] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h191];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h191] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h191];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h192] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h192];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h192] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h192];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h193] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h193];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h193] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h193];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h194] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h194];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h194] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h194];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h195] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h195];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h195] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h195];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h196] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h196];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h196] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h196];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h197] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h197];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h197] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h197];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h198] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h198];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h198] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h198];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h199] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h199];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h199] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h199];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h19f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h19f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h19f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h19f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h1ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h1ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h1ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h1ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h200] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h200];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h200] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h200];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h201] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h201];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h201] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h201];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h202] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h202];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h202] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h202];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h203] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h203];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h203] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h203];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h204] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h204];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h204] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h204];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h205] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h205];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h205] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h205];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h206] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h206];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h206] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h206];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h207] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h207];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h207] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h207];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h208] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h208];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h208] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h208];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h209] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h209];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h209] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h209];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h20f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h20f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h20f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h20f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h210] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h210];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h210] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h210];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h211] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h211];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h211] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h211];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h212] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h212];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h212] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h212];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h213] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h213];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h213] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h213];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h214] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h214];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h214] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h214];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h215] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h215];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h215] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h215];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h216] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h216];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h216] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h216];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h217] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h217];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h217] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h217];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h218] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h218];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h218] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h218];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h219] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h219];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h219] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h219];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h21f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h21f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h21f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h21f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h220] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h220];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h220] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h220];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h221] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h221];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h221] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h221];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h222] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h222];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h222] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h222];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h223] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h223];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h223] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h223];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h224] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h224];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h224] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h224];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h225] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h225];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h225] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h225];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h226] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h226];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h226] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h226];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h227] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h227];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h227] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h227];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h228] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h228];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h228] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h228];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h229] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h229];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h229] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h229];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h22f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h22f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h22f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h22f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h230] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h230];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h230] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h230];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h231] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h231];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h231] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h231];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h232] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h232];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h232] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h232];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h233] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h233];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h233] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h233];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h234] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h234];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h234] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h234];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h235] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h235];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h235] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h235];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h236] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h236];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h236] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h236];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h237] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h237];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h237] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h237];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h238] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h238];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h238] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h238];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h239] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h239];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h239] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h239];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h23f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h23f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h23f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h23f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h240] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h240];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h240] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h240];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h241] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h241];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h241] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h241];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h242] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h242];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h242] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h242];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h243] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h243];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h243] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h243];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h244] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h244];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h244] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h244];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h245] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h245];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h245] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h245];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h246] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h246];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h246] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h246];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h247] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h247];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h247] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h247];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h248] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h248];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h248] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h248];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h249] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h249];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h249] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h249];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h24f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h24f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h24f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h24f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h250] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h250];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h250] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h250];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h251] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h251];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h251] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h251];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h252] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h252];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h252] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h252];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h253] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h253];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h253] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h253];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h254] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h254];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h254] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h254];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h255] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h255];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h255] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h255];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h256] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h256];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h256] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h256];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h257] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h257];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h257] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h257];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h258] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h258];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h258] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h258];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h259] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h259];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h259] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h259];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h25f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h25f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h25f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h25f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h260] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h260];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h260] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h260];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h261] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h261];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h261] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h261];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h262] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h262];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h262] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h262];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h263] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h263];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h263] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h263];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h264] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h264];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h264] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h264];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h265] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h265];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h265] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h265];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h266] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h266];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h266] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h266];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h267] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h267];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h267] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h267];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h268] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h268];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h268] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h268];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h269] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h269];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h269] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h269];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h26f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h26f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h26f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h26f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h270] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h270];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h270] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h270];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h271] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h271];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h271] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h271];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h272] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h272];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h272] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h272];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h273] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h273];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h273] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h273];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h274] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h274];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h274] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h274];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h275] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h275];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h275] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h275];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h276] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h276];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h276] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h276];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h277] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h277];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h277] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h277];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h278] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h278];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h278] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h278];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h279] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h279];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h279] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h279];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h27f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h27f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h27f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h27f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h280] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h280];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h280] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h280];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h281] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h281];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h281] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h281];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h282] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h282];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h282] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h282];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h283] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h283];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h283] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h283];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h284] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h284];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h284] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h284];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h285] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h285];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h285] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h285];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h286] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h286];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h286] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h286];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h287] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h287];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h287] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h287];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h288] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h288];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h288] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h288];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h289] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h289];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h289] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h289];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h28f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h28f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h28f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h28f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h290] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h290];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h290] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h290];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h291] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h291];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h291] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h291];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h292] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h292];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h292] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h292];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h293] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h293];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h293] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h293];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h294] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h294];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h294] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h294];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h295] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h295];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h295] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h295];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h296] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h296];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h296] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h296];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h297] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h297];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h297] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h297];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h298] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h298];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h298] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h298];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h299] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h299];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h299] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h299];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h29f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h29f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h29f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h29f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h2ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h2ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h2ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h2ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h300] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h300];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h300] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h300];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h301] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h301];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h301] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h301];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h302] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h302];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h302] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h302];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h303] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h303];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h303] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h303];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h304] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h304];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h304] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h304];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h305] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h305];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h305] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h305];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h306] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h306];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h306] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h306];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h307] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h307];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h307] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h307];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h308] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h308];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h308] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h308];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h309] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h309];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h309] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h309];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h30f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h30f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h30f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h30f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h310] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h310];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h310] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h310];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h311] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h311];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h311] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h311];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h312] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h312];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h312] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h312];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h313] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h313];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h313] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h313];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h314] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h314];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h314] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h314];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h315] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h315];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h315] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h315];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h316] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h316];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h316] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h316];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h317] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h317];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h317] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h317];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h318] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h318];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h318] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h318];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h319] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h319];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h319] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h319];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h31f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h31f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h31f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h31f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h320] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h320];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h320] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h320];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h321] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h321];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h321] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h321];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h322] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h322];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h322] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h322];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h323] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h323];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h323] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h323];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h324] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h324];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h324] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h324];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h325] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h325];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h325] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h325];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h326] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h326];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h326] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h326];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h327] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h327];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h327] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h327];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h328] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h328];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h328] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h328];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h329] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h329];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h329] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h329];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h32f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h32f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h32f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h32f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h330] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h330];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h330] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h330];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h331] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h331];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h331] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h331];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h332] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h332];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h332] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h332];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h333] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h333];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h333] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h333];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h334] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h334];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h334] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h334];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h335] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h335];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h335] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h335];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h336] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h336];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h336] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h336];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h337] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h337];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h337] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h337];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h338] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h338];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h338] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h338];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h339] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h339];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h339] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h339];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h33f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h33f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h33f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h33f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h340] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h340];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h340] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h340];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h341] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h341];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h341] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h341];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h342] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h342];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h342] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h342];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h343] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h343];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h343] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h343];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h344] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h344];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h344] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h344];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h345] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h345];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h345] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h345];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h346] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h346];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h346] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h346];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h347] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h347];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h347] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h347];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h348] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h348];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h348] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h348];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h349] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h349];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h349] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h349];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h34f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h34f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h34f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h34f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h350] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h350];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h350] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h350];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h351] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h351];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h351] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h351];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h352] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h352];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h352] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h352];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h353] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h353];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h353] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h353];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h354] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h354];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h354] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h354];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h355] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h355];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h355] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h355];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h356] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h356];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h356] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h356];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h357] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h357];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h357] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h357];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h358] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h358];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h358] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h358];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h359] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h359];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h359] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h359];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h35f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h35f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h35f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h35f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h360] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h360];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h360] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h360];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h361] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h361];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h361] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h361];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h362] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h362];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h362] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h362];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h363] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h363];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h363] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h363];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h364] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h364];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h364] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h364];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h365] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h365];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h365] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h365];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h366] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h366];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h366] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h366];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h367] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h367];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h367] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h367];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h368] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h368];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h368] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h368];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h369] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h369];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h369] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h369];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h36f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h36f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h36f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h36f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h370] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h370];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h370] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h370];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h371] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h371];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h371] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h371];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h372] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h372];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h372] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h372];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h373] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h373];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h373] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h373];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h374] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h374];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h374] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h374];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h375] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h375];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h375] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h375];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h376] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h376];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h376] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h376];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h377] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h377];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h377] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h377];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h378] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h378];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h378] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h378];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h379] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h379];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h379] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h379];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h37f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h37f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h37f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h37f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h380] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h380];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h380] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h380];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h381] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h381];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h381] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h381];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h382] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h382];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h382] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h382];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h383] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h383];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h383] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h383];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h384] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h384];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h384] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h384];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h385] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h385];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h385] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h385];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h386] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h386];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h386] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h386];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h387] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h387];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h387] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h387];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h388] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h388];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h388] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h388];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h389] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h389];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h389] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h389];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h38f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h38f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h38f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h38f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h390] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h390];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h390] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h390];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h391] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h391];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h391] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h391];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h392] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h392];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h392] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h392];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h393] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h393];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h393] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h393];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h394] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h394];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h394] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h394];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h395] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h395];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h395] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h395];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h396] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h396];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h396] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h396];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h397] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h397];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h397] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h397];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h398] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h398];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h398] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h398];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h399] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h399];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h399] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h399];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39a] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39a];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39b] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39b];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39c] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39c];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39d] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39d];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39e] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39e];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h39f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h39f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h39f] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h39f];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3a9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3a9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3aa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3aa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ab] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ab];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ac] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ac];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ad] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ad];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ae] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ae];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3af] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3af];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3b9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3b9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ba] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ba];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3be] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3be];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3bf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3bf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3c9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3c9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ca] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ca];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ce] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ce];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3cf] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3cf];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3d9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3d9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3da] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3da];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3db] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3db];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3dc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3dc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3dd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3dd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3de] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3de];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3df] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3df];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3e9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3e9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ea] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ea];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3eb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3eb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ec] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ec];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ed] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ed];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ee] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ee];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ef] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ef];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f0] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f0];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f1] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f1];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f2] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f2];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f3] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f3];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f4] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f4];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f5] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f5];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f6] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f6];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f7] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f7];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f8] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f8];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3f9] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3f9];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fa] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fa];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fb] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fb];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fc] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fc];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fd] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fd];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3fe] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3fe];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[10'h3ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP__[10'h3ff];
    axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[10'h3ff] <= axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD__[10'h3ff];
    array_pointer_delay_0 <= axis_fifo_inst__DOT__wr_addr_reg[32'h9:32'h0];
    if (~(axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[array_pointer_delay_0] | axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[array_pointer_delay_0]) & axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[array_pointer_delay_0]) $display("[%0t] %%loss: axis_fifo_wrapper.axis_fifo_inst__DOT__mem 'd31 'd0 axis_fifo_wrapper.array_pointer_delay_0 PartSelect ptr=h%h", $time , array_pointer_delay_0) /*debug_display_flowguard*/; 
  end

  always @(posedge clk) begin
    if (rst) TASKPASS_cycle_counter <= 64'h0; 
    else TASKPASS_cycle_counter <= (TASKPASS_cycle_counter + 64'h1);
  end
  wire display_cond_0 ;
  assign display_cond_0 = (axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____ASSIGN_Q__ && !axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____GOOD_Q__ && !axis_fifo_inst__DOT__mem_read_data_reg__BRA__31__03A0__KET____PROP_Q__);
  wire display_cond_1 ;
  assign display_cond_1 = (axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____ASSIGN_Q__[array_pointer_delay_0] && !axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____GOOD_Q__[array_pointer_delay_0] && !axis_fifo_inst__DOT__mem__BRA__31__03A0__KET____PROP_Q__[array_pointer_delay_0]);

  ila_losscheck
  ila_inst_0
  (
    .clk(clk),
    .probe0({ display_cond_0, display_cond_1, TASKPASS_cycle_counter, array_pointer_delay_0 }),
    .probe1(display_cond_0 || display_cond_1)
  );


endmodule
