`define HLS_NAME mobilenet
