`define HLS_NAME top
