`define HLS_NAME rendering
