`define HLS_NAME optical_flow
