`include "cl_fpgarr_defs.svh"
////////////////////////////////////////////////////////////////////////////
// axi interconnect for merging CL pcim requests with the pcim requests
// converted from interrupt
// This is just a workaround to support interrupt in the happen-before trace
////////////////////////////////////////////////////////////////////////////
module rr_cl_irq2pcim_interconnect (
  input wire clk,
  input wire rstn,
  rr_axi_bus_t.master rr_pcim_bus,
  rr_axi_bus_t.master irq_pcim_bus,
  rr_axi_bus_t.slave rr_irq_pcim_bus
);
localparam int NUM_SLV = 2;
if (CL_PCIM_AXI_ID_WIDTH + $clog2(NUM_SLV) > PCIM_INTERCONNECT_AXI_ID_WIDTH)
  $error("AXI ID allocation is invalid: irq_pcim NUM_SLV %d, CL_PCIM_AXI_ID_WIDTH %d, PCIM_INTERCONNECT_AXI_ID_WIDTH %d",
    NUM_SLV, CL_PCIM_AXI_ID_WIDTH, PCIM_INTERCONNECT_AXI_ID_WIDTH);
// NOTE: S00 is READ WRITE, for rr_pcim
//       S01 is WRITE ONLY, for irq_pcim
rr_irq_pcim_interconnect irq_pcim_interconnect_inst (
  .ACLK(clk),
  .ARESETN(rstn),
  /* the single output master bus connecting to the pcim_axi_interconnect */
  .M00_AXI_araddr(rr_irq_pcim_bus.araddr),
  .M00_AXI_arburst(),
  .M00_AXI_arcache(),
  .M00_AXI_arid(rr_irq_pcim_bus.arid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
  .M00_AXI_arlen(rr_irq_pcim_bus.arlen),
  .M00_AXI_arlock(),
  .M00_AXI_arprot(),
  .M00_AXI_arqos(),
  .M00_AXI_arready(rr_irq_pcim_bus.arready),
  .M00_AXI_arregion(),
  .M00_AXI_arsize(rr_irq_pcim_bus.arsize),
  .M00_AXI_arvalid(rr_irq_pcim_bus.arvalid),
  .M00_AXI_awaddr(rr_irq_pcim_bus.awaddr),
  .M00_AXI_awburst(),
  .M00_AXI_awcache(),
  .M00_AXI_awid(rr_irq_pcim_bus.awid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
  .M00_AXI_awlen(rr_irq_pcim_bus.awlen),
  .M00_AXI_awlock(),
  .M00_AXI_awprot(),
  .M00_AXI_awqos(),
  .M00_AXI_awready(rr_irq_pcim_bus.awready),
  .M00_AXI_awregion(),
  .M00_AXI_awsize(rr_irq_pcim_bus.awsize),
  .M00_AXI_awvalid(rr_irq_pcim_bus.awvalid),
  .M00_AXI_bid(rr_irq_pcim_bus.bid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
  .M00_AXI_bready(rr_irq_pcim_bus.bready),
  .M00_AXI_bresp(rr_irq_pcim_bus.bresp),
  .M00_AXI_bvalid(rr_irq_pcim_bus.bvalid),
  .M00_AXI_rdata(rr_irq_pcim_bus.rdata),
  .M00_AXI_rid(rr_irq_pcim_bus.rid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
  .M00_AXI_rlast(rr_irq_pcim_bus.rlast),
  .M00_AXI_rready(rr_irq_pcim_bus.rready),
  .M00_AXI_rresp(rr_irq_pcim_bus.rresp),
  .M00_AXI_rvalid(rr_irq_pcim_bus.rvalid),
  .M00_AXI_wdata(rr_irq_pcim_bus.wdata),
  .M00_AXI_wlast(rr_irq_pcim_bus.wlast),
  .M00_AXI_wready(rr_irq_pcim_bus.wready),
  .M00_AXI_wstrb(rr_irq_pcim_bus.wstrb),
  .M00_AXI_wvalid(rr_irq_pcim_bus.wvalid),
  /* cl pcim requests (READ WRITE) */
  .S00_AXI_araddr(rr_pcim_bus.araddr),
  .S00_AXI_arburst(2'b1), // INCR
  .S00_AXI_arcache(4'b00),
  .S00_AXI_arid(rr_pcim_bus.arid[CL_PCIM_AXI_ID_WIDTH-1:0]),
  .S00_AXI_arlen(rr_pcim_bus.arlen),
  .S00_AXI_arlock(1'b0),
  .S00_AXI_arprot(3'b00),
  .S00_AXI_arqos(4'b0),
  .S00_AXI_arready(rr_pcim_bus.arready),
  .S00_AXI_arregion(4'b0),
  .S00_AXI_arsize(rr_pcim_bus.arsize),
  .S00_AXI_arvalid(rr_pcim_bus.arvalid),
  .S00_AXI_awaddr(rr_pcim_bus.awaddr),
  .S00_AXI_awburst(2'b1),
  .S00_AXI_awcache(4'b00),
  .S00_AXI_awid(rr_pcim_bus.awid[CL_PCIM_AXI_ID_WIDTH-1:0]),
  .S00_AXI_awlen(rr_pcim_bus.awlen),
  .S00_AXI_awlock(1'b0),
  .S00_AXI_awprot(3'b00),
  .S00_AXI_awqos(4'b0),
  .S00_AXI_awready(rr_pcim_bus.awready),
  .S00_AXI_awregion(4'b0),
  .S00_AXI_awsize(rr_pcim_bus.awsize),
  .S00_AXI_awvalid(rr_pcim_bus.awvalid),
  .S00_AXI_bid(rr_pcim_bus.bid[CL_PCIM_AXI_ID_WIDTH-1:0]),
  .S00_AXI_bready(rr_pcim_bus.bready),
  .S00_AXI_bresp(rr_pcim_bus.bresp),
  .S00_AXI_bvalid(rr_pcim_bus.bvalid),
  .S00_AXI_rdata(rr_pcim_bus.rdata),
  .S00_AXI_rid(rr_pcim_bus.rid[CL_PCIM_AXI_ID_WIDTH-1:0]),
  .S00_AXI_rlast(rr_pcim_bus.rlast),
  .S00_AXI_rready(rr_pcim_bus.rready),
  .S00_AXI_rresp(rr_pcim_bus.rresp),
  .S00_AXI_rvalid(rr_pcim_bus.rvalid),
  .S00_AXI_wdata(rr_pcim_bus.wdata),
  .S00_AXI_wlast(rr_pcim_bus.wlast),
  .S00_AXI_wready(rr_pcim_bus.wready),
  .S00_AXI_wstrb(rr_pcim_bus.wstrb),
  .S00_AXI_wvalid(rr_pcim_bus.wvalid),
  /* interrupt requests => pcim requests (WRITE ONLY) */
  .S01_AXI_awaddr(irq_pcim_bus.awaddr),
  .S01_AXI_awburst(2'b1),
  .S01_AXI_awcache(4'b00),
  .S01_AXI_awid(irq_pcim_bus.awid[CL_PCIM_AXI_ID_WIDTH-1:0]),
  .S01_AXI_awlen(irq_pcim_bus.awlen),
  .S01_AXI_awlock(1'b0),
  .S01_AXI_awprot(3'b00),
  .S01_AXI_awqos(4'b0),
  .S01_AXI_awready(irq_pcim_bus.awready),
  .S01_AXI_awregion(4'b0),
  .S01_AXI_awsize(irq_pcim_bus.awsize),
  .S01_AXI_awvalid(irq_pcim_bus.awvalid),
  .S01_AXI_bid(irq_pcim_bus.bid[CL_PCIM_AXI_ID_WIDTH-1:0]),
  .S01_AXI_bready(irq_pcim_bus.bready),
  .S01_AXI_bresp(irq_pcim_bus.bresp),
  .S01_AXI_bvalid(irq_pcim_bus.bvalid),
  .S01_AXI_wdata(irq_pcim_bus.wdata),
  .S01_AXI_wlast(irq_pcim_bus.wlast),
  .S01_AXI_wready(irq_pcim_bus.wready),
  .S01_AXI_wstrb(irq_pcim_bus.wstrb),
  .S01_AXI_wvalid(irq_pcim_bus.wvalid)
);
endmodule
