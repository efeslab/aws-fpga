`define HLS_NAME nbody
