`define HLS_NAME calc_0
