`define HLS_NAME bellman_ford
