`define HLS_NAME hashing_kernel
