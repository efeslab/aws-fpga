module axil_rr_mstr (
   input clk,
   input sync_rst_n,
   axi_lite_bus_t.to_master axil_in,
   
   axi_lite_bus_t.to_slave axil_out,
);

axi
endmodule
