`include "cl_fpgarr_defs.svh"
////////////////////////////////////////////////////////////////////////////
// axi interconnect for sharing single shell pcim bus across the logging
// writeback module and the user pcim bus
////////////////////////////////////////////////////////////////////////////
module rr_storage_pcim_axi_interconnect (
   input wire clk,
   input wire rstn,
   rr_axi_bus_t.master logging_wb_bus,
   rr_axi_bus_t.master validation_wb_bus,
   rr_axi_bus_t.master cl_pcim_bus,
   rr_axi_bus_t.slave sh_pcim_bus
);

localparam int AXI_ID_WIDTH = 16;
localparam int NUM_SLV = 3;
if (PCIM_INTERCONNECT_AXI_ID_WIDTH + $clog2(NUM_SLV) > AXI_ID_WIDTH)
   $error("ID allocation is invalid: NUM_SLV %d, PCIM_INTERCONNECT_AXI_ID_WIDTH %d",
      NUM_SLV, PCIM_INTERCONNECT_AXI_ID_WIDTH);
// TODO: is this dont_touch necessary?
// NOTE: S00 is READ WRITE
//       S01 is WRITE ONLY
//       S02 is READ WRITE
(* dont_touch = "true" *) rr_pcim_axi_interconnect pcim_interconnect_inst (
   .ACLK(clk),
   .ARESETN(rstn),
   /* the single output master bus connecting to the shell*/
   .M00_AXI_araddr(sh_pcim_bus.araddr),
   .M00_AXI_arburst(),
   .M00_AXI_arcache(),
   .M00_AXI_arid(sh_pcim_bus.arid),
   .M00_AXI_arlen(sh_pcim_bus.arlen),
   .M00_AXI_arlock(),
   .M00_AXI_arprot(),
   .M00_AXI_arqos(),
   .M00_AXI_arready(sh_pcim_bus.arready),
   .M00_AXI_arregion(),
   .M00_AXI_arsize(sh_pcim_bus.arsize),
   .M00_AXI_arvalid(sh_pcim_bus.arvalid),
   .M00_AXI_awaddr(sh_pcim_bus.awaddr),
   .M00_AXI_awburst(),
   .M00_AXI_awcache(),
   .M00_AXI_awid(sh_pcim_bus.awid),
   .M00_AXI_awlen(sh_pcim_bus.awlen),
   .M00_AXI_awlock(),
   .M00_AXI_awprot(),
   .M00_AXI_awqos(),
   .M00_AXI_awready(sh_pcim_bus.awready),
   .M00_AXI_awregion(),
   .M00_AXI_awsize(sh_pcim_bus.awsize),
   .M00_AXI_awvalid(sh_pcim_bus.awvalid),
   .M00_AXI_bid(sh_pcim_bus.bid),
   .M00_AXI_bready(sh_pcim_bus.bready),
   .M00_AXI_bresp(sh_pcim_bus.bresp),
   .M00_AXI_bvalid(sh_pcim_bus.bvalid),
   .M00_AXI_rdata(sh_pcim_bus.rdata),
   .M00_AXI_rid(sh_pcim_bus.rid),
   .M00_AXI_rlast(sh_pcim_bus.rlast),
   .M00_AXI_rready(sh_pcim_bus.rready),
   .M00_AXI_rresp(sh_pcim_bus.rresp),
   .M00_AXI_rvalid(sh_pcim_bus.rvalid),
   .M00_AXI_wdata(sh_pcim_bus.wdata),
   .M00_AXI_wlast(sh_pcim_bus.wlast),
   .M00_AXI_wready(sh_pcim_bus.wready),
   .M00_AXI_wstrb(sh_pcim_bus.wstrb),
   .M00_AXI_wvalid(sh_pcim_bus.wvalid),
   /* logging writeback bus (generated by fpgarr for record/replay) */
   .S00_AXI_araddr(logging_wb_bus.araddr),
   .S00_AXI_arburst(2'b1), // INCR
   .S00_AXI_arcache(4'b00),
   .S00_AXI_arid(logging_wb_bus.arid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S00_AXI_arlen(logging_wb_bus.arlen),
   .S00_AXI_arlock(1'b0),
   .S00_AXI_arprot(3'b00),
   .S00_AXI_arqos(4'b0),
   .S00_AXI_arready(logging_wb_bus.arready),
   .S00_AXI_arregion(4'b0),
   .S00_AXI_arsize(logging_wb_bus.arsize),
   .S00_AXI_arvalid(logging_wb_bus.arvalid),
   .S00_AXI_awaddr(logging_wb_bus.awaddr),
   .S00_AXI_awburst(2'b1),
   .S00_AXI_awcache(4'b00),
   .S00_AXI_awid(logging_wb_bus.awid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S00_AXI_awlen(logging_wb_bus.awlen),
   .S00_AXI_awlock(1'b0),
   .S00_AXI_awprot(3'b00),
   .S00_AXI_awqos(4'b0),
   .S00_AXI_awready(logging_wb_bus.awready),
   .S00_AXI_awregion(4'b0),
   .S00_AXI_awsize(logging_wb_bus.awsize),
   .S00_AXI_awvalid(logging_wb_bus.awvalid),
   .S00_AXI_bid(logging_wb_bus.bid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S00_AXI_bready(logging_wb_bus.bready),
   .S00_AXI_bresp(logging_wb_bus.bresp),
   .S00_AXI_bvalid(logging_wb_bus.bvalid),
   .S00_AXI_rdata(logging_wb_bus.rdata),
   .S00_AXI_rid(logging_wb_bus.rid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S00_AXI_rlast(logging_wb_bus.rlast),
   .S00_AXI_rready(logging_wb_bus.rready),
   .S00_AXI_rresp(logging_wb_bus.rresp),
   .S00_AXI_rvalid(logging_wb_bus.rvalid),
   .S00_AXI_wdata(logging_wb_bus.wdata),
   .S00_AXI_wlast(logging_wb_bus.wlast),
   .S00_AXI_wready(logging_wb_bus.wready),
   .S00_AXI_wstrb(logging_wb_bus.wstrb),
   .S00_AXI_wvalid(logging_wb_bus.wvalid),
   /* validation writeback bus (generated by fpgarr for output validation) */
   .S01_AXI_araddr(64'b0),
   .S01_AXI_arburst(2'b1),
   .S01_AXI_arcache(4'b00),
   .S01_AXI_arid(14'b0),
   .S01_AXI_arlen(8'b0),
   .S01_AXI_arlock(1'b0),
   .S01_AXI_arprot(3'b00),
   .S01_AXI_arqos(4'b0),
   .S01_AXI_arready(),
   .S01_AXI_arregion(4'b0),
   .S01_AXI_arsize(3'b0),
   .S01_AXI_arvalid(1'b0),
   .S01_AXI_awaddr(validation_wb_bus.awaddr),
   .S01_AXI_awburst(2'b1),
   .S01_AXI_awcache(4'b00),
   .S01_AXI_awid(validation_wb_bus.awid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S01_AXI_awlen(validation_wb_bus.awlen),
   .S01_AXI_awlock(1'b0),
   .S01_AXI_awprot(3'b00),
   .S01_AXI_awqos(4'b0),
   .S01_AXI_awready(validation_wb_bus.awready),
   .S01_AXI_awregion(4'b0),
   .S01_AXI_awsize(validation_wb_bus.awsize),
   .S01_AXI_awvalid(validation_wb_bus.awvalid),
   .S01_AXI_bid(validation_wb_bus.bid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S01_AXI_bready(validation_wb_bus.bready),
   .S01_AXI_bresp(validation_wb_bus.bresp),
   .S01_AXI_bvalid(validation_wb_bus.bvalid),
   .S01_AXI_rdata(),
   .S01_AXI_rid(),
   .S01_AXI_rlast(),
   .S01_AXI_rready(1'b1),
   .S01_AXI_rresp(),
   .S01_AXI_rvalid(),
   .S01_AXI_wdata(validation_wb_bus.wdata),
   .S01_AXI_wlast(validation_wb_bus.wlast),
   .S01_AXI_wready(validation_wb_bus.wready),
   .S01_AXI_wstrb(validation_wb_bus.wstrb),
   .S01_AXI_wvalid(validation_wb_bus.wvalid),
   /* cl pcim bus (should be taken care of in rr) */
   .S02_AXI_araddr(cl_pcim_bus.araddr),
   .S02_AXI_arburst(2'b1), // INCR
   .S02_AXI_arcache(4'b00),
   .S02_AXI_arid(cl_pcim_bus.arid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S02_AXI_arlen(cl_pcim_bus.arlen),
   .S02_AXI_arlock(1'b0),
   .S02_AXI_arprot(3'b00),
   .S02_AXI_arqos(4'b0),
   .S02_AXI_arready(cl_pcim_bus.arready),
   .S02_AXI_arregion(4'b0),
   .S02_AXI_arsize(cl_pcim_bus.arsize),
   .S02_AXI_arvalid(cl_pcim_bus.arvalid),
   .S02_AXI_awaddr(cl_pcim_bus.awaddr),
   .S02_AXI_awburst(2'b1),
   .S02_AXI_awcache(4'b00),
   .S02_AXI_awid(cl_pcim_bus.awid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S02_AXI_awlen(cl_pcim_bus.awlen),
   .S02_AXI_awlock(1'b0),
   .S02_AXI_awprot(3'b00),
   .S02_AXI_awqos(4'b0),
   .S02_AXI_awready(cl_pcim_bus.awready),
   .S02_AXI_awregion(4'b0),
   .S02_AXI_awsize(cl_pcim_bus.awsize),
   .S02_AXI_awvalid(cl_pcim_bus.awvalid),
   .S02_AXI_bid(cl_pcim_bus.bid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S02_AXI_bready(cl_pcim_bus.bready),
   .S02_AXI_bresp(cl_pcim_bus.bresp),
   .S02_AXI_bvalid(cl_pcim_bus.bvalid),
   .S02_AXI_rdata(cl_pcim_bus.rdata),
   .S02_AXI_rid(cl_pcim_bus.rid[PCIM_INTERCONNECT_AXI_ID_WIDTH-1:0]),
   .S02_AXI_rlast(cl_pcim_bus.rlast),
   .S02_AXI_rready(cl_pcim_bus.rready),
   .S02_AXI_rresp(cl_pcim_bus.rresp),
   .S02_AXI_rvalid(cl_pcim_bus.rvalid),
   .S02_AXI_wdata(cl_pcim_bus.wdata),
   .S02_AXI_wlast(cl_pcim_bus.wlast),
   .S02_AXI_wready(cl_pcim_bus.wready),
   .S02_AXI_wstrb(cl_pcim_bus.wstrb),
   .S02_AXI_wvalid(cl_pcim_bus.wvalid)
);

// mask the read interface of the validation_wb_bus (since it is write-only)
assign validation_wb_bus.arready = 1;
assign validation_wb_bus.rvalid = 0;
// clear the higher reserved id for all slaves
`define CLEAR_PCIM_AXI_ID(bus) \
   assign bus.bid[AXI_ID_WIDTH-1:PCIM_INTERCONNECT_AXI_ID_WIDTH] = 0; \
   assign bus.rid[AXI_ID_WIDTH-1:PCIM_INTERCONNECT_AXI_ID_WIDTH] = 0
`CLEAR_PCIM_AXI_ID(logging_wb_bus);
`CLEAR_PCIM_AXI_ID(validation_wb_bus);
`CLEAR_PCIM_AXI_ID(cl_pcim_bus);

`ifdef DEBUG_INTERCONNECT
pcim_dbg_cnt dbg_record_cnt (
   .clk(clk), .rstn(rstn),
   .bus(logging_wb_bus)
);
pcim_dbg_cnt dbg_validate_cnt (
   .clk(clk), .rstn(rstn),
   .bus(validation_wb_bus)
);
pcim_dbg_cnt dbg_cl_cnt (
   .clk(clk), .rstn(rstn),
   .bus(cl_pcim_bus)
);
pcim_dbg_cnt dbg_sh_cnt (
   .clk(clk), .rstn(rstn),
   .bus(sh_pcim_bus)
);
`endif
endmodule
