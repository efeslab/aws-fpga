`define HLS_NAME SgdLR
