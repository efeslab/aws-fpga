module rr_packed2writeback_bus (
   input wire clk,
   input wire rstn,
   rr_packed_logging_bus_t.C in,
   rr_stream_bus_t.P out
);

// parameter check
generate
   if (in.LOGB_CHANNEL_CNT + in.LOGE_CHANNEL_CNT + in.FULL_WIDTH
       != out.FULL_WIDTH)
    $error("Writeback FULL_WIDTH mismatch: logb W%d, loge W%d, packed_logb_data W%d, writeback W%d\n",
      in.LOGB_CHANNEL_CNT, in.LOGE_CHANNEL_CNT, in.FULL_WIDTH, out.FULL_WIDTH);
endgenerate

// loge_valid_output is the signal outputting to the writeback_bus
// loge_valid_output[i] shows whether one (and can only be one) transaction has
// finished on channel[i] between now (some logb_valid are true) and the last
// time some logb are valid.
// if logb_valid[i] && loge_valid[i], which only happen if the transaction
// really lasts for only one cycle (ready was asserted in advance)
logic [in.LOGE_CHANNEL_CNT-1:0] loge_valid_out;

assign out.valid = in.plogb.any_valid;
assign in.ready = out.ready;
assign out.len = out.valid?
   (in.plogb.len + out.OFFSET_WIDTH'(in.LOGB_CHANNEL_CNT + in.LOGE_CHANNEL_CNT))
   : 0;
// from LSB to MSB:
// logb_valid, loge_valid, packed_logb_data
assign out.data = {in.plogb.data, loge_valid_out, in.logb_valid};

// buf loge_valid if there is no valid logb to send
always @(posedge clk)
if (!rstn)
   loge_valid_out <= 0;
else
   for (int i=0; i < in.LOGE_CHANNEL_CNT; i=i+1)
      if (out.valid && in.loge_valid[i])
         loge_valid_out[i] <= 1;
      else if (out.valid && !in.loge_valid[i])
         loge_valid_out[i] <= 0;
      else if (!out.valid && in.loge_valid[i]) begin
         loge_valid_out[i] <= 1;
         no_loge_overwrite: assert(!loge_valid_out[i]);
      end
      else // !out.valid && !in.loge_valid[i]
         loge_valid_out[i] <= loge_valid_out[i];
endmodule

////////////////////////////////////////////////////////////////////////////
// axi interconnect for sharing single shell pcim bus across the logging
// writeback module and the user pcim bus
////////////////////////////////////////////////////////////////////////////
module rr_storage_pcim_axi_interconnect (
   input wire clk,
   input wire rstn,
   rr_axi_bus_t.master logging_wb_bus,
   rr_axi_bus_t.master cl_pcim_bus,
   rr_axi_bus_t.slave sh_pcim_bus
);

rr_pcim_axi_interconnect pcim_interconnect_inst (
   .ACLK(clk),
   .ARESETN(rstn),
   /* the single output master bus connecting to the shell*/
   .M00_AXI_araddr(sh_pcim_bus.araddr),
   .M00_AXI_arburst(),
   .M00_AXI_arcache(),
   .M00_AXI_arid(sh_pcim_bus.arid),
   .M00_AXI_arlen(sh_pcim_bus.arlen),
   .M00_AXI_arlock(),
   .M00_AXI_arprot(),
   .M00_AXI_arqos(),
   .M00_AXI_arready(sh_pcim_bus.arready),
   .M00_AXI_arregion(),
   .M00_AXI_arsize(sh_pcim_bus.arsize),
   .M00_AXI_arvalid(sh_pcim_bus.arvalid),
   .M00_AXI_awaddr(sh_pcim_bus.awaddr),
   .M00_AXI_awburst(),
   .M00_AXI_awcache(),
   .M00_AXI_awid(sh_pcim_bus.awid),
   .M00_AXI_awlen(sh_pcim_bus.awlen),
   .M00_AXI_awlock(),
   .M00_AXI_awprot(),
   .M00_AXI_awqos(),
   .M00_AXI_awready(sh_pcim_bus.awready),
   .M00_AXI_awregion(),
   .M00_AXI_awsize(sh_pcim_bus.awsize),
   .M00_AXI_awvalid(sh_pcim_bus.awvalid),
   .M00_AXI_bid(sh_pcim_bus.bid),
   .M00_AXI_bready(sh_pcim_bus.bready),
   .M00_AXI_bresp(sh_pcim_bus.bresp),
   .M00_AXI_bvalid(sh_pcim_bus.bvalid),
   .M00_AXI_rdata(sh_pcim_bus.rdata),
   .M00_AXI_rid(sh_pcim_bus.rid),
   .M00_AXI_rlast(sh_pcim_bus.rlast),
   .M00_AXI_rready(sh_pcim_bus.rready),
   .M00_AXI_rresp(sh_pcim_bus.rresp),
   .M00_AXI_rvalid(sh_pcim_bus.rvalid),
   .M00_AXI_wdata(sh_pcim_bus.wdata),
   .M00_AXI_wlast(sh_pcim_bus.wlast),
   .M00_AXI_wready(sh_pcim_bus.wready),
   .M00_AXI_wstrb(sh_pcim_bus.wstrb),
   .M00_AXI_wvalid(sh_pcim_bus.wvalid),
   /* logging writeback bus (generated by rr) */
   .S00_AXI_araddr(logging_wb_bus.araddr),
   .S00_AXI_arburst(2'b1), // INCR
   .S00_AXI_arcache(4'b00),
   .S00_AXI_arid(logging_wb_bus.arid[14:0]),
   .S00_AXI_arlen(logging_wb_bus.arlen),
   .S00_AXI_arlock(1'b0),
   .S00_AXI_arprot(3'b00),
   .S00_AXI_arqos(4'b0),
   .S00_AXI_arready(logging_wb_bus.arready),
   .S00_AXI_arregion(4'b0),
   .S00_AXI_arsize(logging_wb_bus.arsize),
   .S00_AXI_arvalid(logging_wb_bus.arvalid),
   .S00_AXI_awaddr(logging_wb_bus.awaddr),
   .S00_AXI_awburst(2'b1),
   .S00_AXI_awcache(4'b00),
   .S00_AXI_awid(logging_wb_bus.awid[14:0]),
   .S00_AXI_awlen(logging_wb_bus.awlen),
   .S00_AXI_awlock(1'b0),
   .S00_AXI_awprot(3'b00),
   .S00_AXI_awqos(4'b0),
   .S00_AXI_awready(logging_wb_bus.awready),
   .S00_AXI_awregion(4'b0),
   .S00_AXI_awsize(logging_wb_bus.awsize),
   .S00_AXI_awvalid(logging_wb_bus.awvalid),
   .S00_AXI_bid(logging_wb_bus.bid[14:0]),
   .S00_AXI_bready(logging_wb_bus.bready),
   .S00_AXI_bresp(logging_wb_bus.bresp),
   .S00_AXI_bvalid(logging_wb_bus.bvalid),
   .S00_AXI_rdata(logging_wb_bus.rdata),
   .S00_AXI_rid(logging_wb_bus.rid[14:0]),
   .S00_AXI_rlast(logging_wb_bus.rlast),
   .S00_AXI_rready(logging_wb_bus.rready),
   .S00_AXI_rresp(logging_wb_bus.rresp),
   .S00_AXI_rvalid(logging_wb_bus.rvalid),
   .S00_AXI_wdata(logging_wb_bus.wdata),
   .S00_AXI_wlast(logging_wb_bus.wlast),
   .S00_AXI_wready(logging_wb_bus.wready),
   .S00_AXI_wstrb(logging_wb_bus.wstrb),
   .S00_AXI_wvalid(logging_wb_bus.wvalid),
   /* cl pcim bus (should be taken care of in rr) */
   .S01_AXI_araddr(cl_pcim_bus.araddr),
   .S01_AXI_arburst(2'b1), // INCR
   .S01_AXI_arcache(4'b00),
   .S01_AXI_arid(cl_pcim_bus.arid[14:0]),
   .S01_AXI_arlen(cl_pcim_bus.arlen),
   .S01_AXI_arlock(1'b0),
   .S01_AXI_arprot(3'b00),
   .S01_AXI_arqos(4'b0),
   .S01_AXI_arready(cl_pcim_bus.arready),
   .S01_AXI_arregion(4'b0),
   .S01_AXI_arsize(cl_pcim_bus.arsize),
   .S01_AXI_arvalid(cl_pcim_bus.arvalid),
   .S01_AXI_awaddr(cl_pcim_bus.awaddr),
   .S01_AXI_awburst(2'b1),
   .S01_AXI_awcache(4'b00),
   .S01_AXI_awid(cl_pcim_bus.awid[14:0]),
   .S01_AXI_awlen(cl_pcim_bus.awlen),
   .S01_AXI_awlock(1'b0),
   .S01_AXI_awprot(3'b00),
   .S01_AXI_awqos(4'b0),
   .S01_AXI_awready(cl_pcim_bus.awready),
   .S01_AXI_awregion(4'b0),
   .S01_AXI_awsize(cl_pcim_bus.awsize),
   .S01_AXI_awvalid(cl_pcim_bus.awvalid),
   .S01_AXI_bid(cl_pcim_bus.bid[14:0]),
   .S01_AXI_bready(cl_pcim_bus.bready),
   .S01_AXI_bresp(cl_pcim_bus.bresp),
   .S01_AXI_bvalid(cl_pcim_bus.bvalid),
   .S01_AXI_rdata(cl_pcim_bus.rdata),
   .S01_AXI_rid(cl_pcim_bus.rid[14:0]),
   .S01_AXI_rlast(cl_pcim_bus.rlast),
   .S01_AXI_rready(cl_pcim_bus.rready),
   .S01_AXI_rresp(cl_pcim_bus.rresp),
   .S01_AXI_rvalid(cl_pcim_bus.rvalid),
   .S01_AXI_wdata(cl_pcim_bus.wdata),
   .S01_AXI_wlast(cl_pcim_bus.wlast),
   .S01_AXI_wready(cl_pcim_bus.wready),
   .S01_AXI_wstrb(cl_pcim_bus.wstrb),
   .S01_AXI_wvalid(cl_pcim_bus.wvalid)
);
endmodule

/*
 * A better structure in my mind.
 * Summary of the requirement:
 * ===> Variable length input (0..WIDTH)
 *             Fixed 512 output (AXI_WIDTH) ===>
 * A [2*WIDTH-1:0] (shift register?) B
 * Four cases to consider:
 * B_next
 * B
 * 1. !in, !out B_next = B
 * 2. in, !out
 *    B_next[B_len +: WIDTH] = in
 * 3. !in, out
 *    B_next[0 +: WIDTH-AXI_WIDTH] = B[AXI_WIDTH +: WIDTH-AXI_WIDTH]
 *    out[AXI_WIDTH-1:0] = B[0 +: AXI_WIDTH]
 * 4. in, out
 *    B_next[0 +: WIDTH-AXI_WIDTH] = B[AXI_WIDTH +: WIDTH-AXI_WIDTH]
 *    B_next[B_len - AXI_WIDTH +: WIDTH] = in
 *    out[AXI_WIDTH-1:0] = B[0 +: AXI_WIDTH]
 */
module rr_writeback #(
    parameter WIDTH = 2500,
    parameter AXI_WIDTH = 512,
    parameter OFFSETWIDTH = 32,
    parameter AXI_ADDR_WIDTH = 64) (
    input clk,
    input sync_rst_n,
    // cfg_max_payload: see https://github.com/aws/aws-fpga/blob/master/hdk/docs/AWS_Shell_Interface_Specification.md#pcim-interface----axi-4-for-outbound-pcie-transactions-cl-is-master-shell-is-slave-512-bit
    input logic [1:0] cfg_max_payload,

    input logic din_valid,
    output logic din_ready,
    input logic finish,
    input logic [WIDTH-1:0] din,
    input logic [OFFSETWIDTH-1:0] din_width,

    rr_axi_bus_t.slave axi_out,
    input logic [AXI_ADDR_WIDTH-1:0] buf_addr,
    input logic [AXI_ADDR_WIDTH-1:0] buf_size,
    input logic buf_update,

    // When there's a buffer overflow, the interrupt will be triggerred
    output logic interrupt
);

    localparam NSTAGES = (WIDTH - 1) / AXI_WIDTH + 1;
    localparam EXT_WIDTH = NSTAGES * AXI_WIDTH;

    logic [WIDTH-1:0] in_fifo_out;
    logic [EXT_WIDTH-1:0] in_fifo_out_wrap;
    logic [OFFSETWIDTH-1:0] in_fifo_out_width;
    logic in_fifo_rd_en;
    logic in_fifo_full, in_fifo_almfull, in_fifo_empty;

    assign in_fifo_out_wrap = EXT_WIDTH'(in_fifo_out);

    merged_fifo #(
        .WIDTH(WIDTH+OFFSETWIDTH),
        .ALMFULL_THRESHOLD(12))
    mfifo_inst_in(
        .clk(clk),
        .rst(~sync_rst_n),
        .din({din,din_width}),
        .dout({in_fifo_out,in_fifo_out_width}),
        .wr_en(din_valid),
        .rd_en(in_fifo_rd_en),
        .full(in_fifo_full),
        .almfull(in_fifo_almfull),
        .empty(in_fifo_empty)
    );

    logic [AXI_WIDTH-1:0] out_fifo_out, out_fifo_in, out_fifo_in_q, out_fifo_in_qq;
    logic out_fifo_rd_en, out_fifo_wr_en, out_fifo_wr_en_q, out_fifo_wr_en_qq;
    logic out_fifo_full, out_fifo_almfull, out_fifo_empty;

    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            out_fifo_wr_en_qq <= 0;
        end else begin
            out_fifo_in_q <= out_fifo_in;
            out_fifo_in_qq <= out_fifo_in_q;
            out_fifo_wr_en_q <= out_fifo_wr_en;
            out_fifo_wr_en_qq <= out_fifo_wr_en_q;
        end
    end

    merged_fifo #(
        .WIDTH(AXI_WIDTH),
        .ALMFULL_THRESHOLD(12))
    mfifo_inst_out(
        .clk(clk),
        .rst(~sync_rst_n),
        .din(out_fifo_in_qq),
        .dout(out_fifo_out),
        .wr_en(out_fifo_wr_en_qq),
        .rd_en(out_fifo_rd_en),
        .full(out_fifo_full),
        .almfull(out_fifo_almfull),
        .empty(out_fifo_empty)
    );

    logic [OFFSETWIDTH-1:0] unhandled_size;
    logic [AXI_WIDTH-1:0] unhandled [NSTAGES-1:0];
    logic [AXI_WIDTH-1:0] leftover;
    logic [$clog2(AXI_WIDTH):0] leftover_size;
    logic [$clog2(NSTAGES):0] curr;
    logic do_finish;

    assign in_fifo_rd_en = ~in_fifo_empty && ~out_fifo_almfull && unhandled_size <= AXI_WIDTH;

    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            unhandled_size <= 0;
            leftover_size <= 0;
            curr <= 0;
            do_finish <= 0;
            out_fifo_in <= 0;
        end else begin
            if (finish) begin
                do_finish <= 1;
            end

            if (in_fifo_rd_en) begin
                curr <= 0;
                unhandled_size <= in_fifo_out_width;
                for (int i = 0; i < NSTAGES; i++) begin
                    unhandled[i] <= in_fifo_out_wrap[i*AXI_WIDTH+:AXI_WIDTH];
                end
            end else if (curr + 1 <= NSTAGES) begin
                curr <= curr + 1;
                if (unhandled_size >= AXI_WIDTH) begin
                    unhandled_size <= unhandled_size - AXI_WIDTH;
                end else begin
                    unhandled_size <= 0;
                end
            end

`ifdef TEST_DIRECT_CONNECT
            if (unhandled_size >= 0) begin
                out_fifo_in <= unhandled[curr];
                out_fifo_wr_en <= 1;
            end else begin
                out_fifo_wr_en <= 0;
            end
`else
            if (unhandled_size >= AXI_WIDTH) begin
                leftover_size <= leftover_size;
                leftover <= unhandled[curr] >> (AXI_WIDTH - leftover_size);
                out_fifo_in <= (unhandled[curr] << leftover_size) | (leftover & (AXI_WIDTH'(-1) >> (AXI_WIDTH - leftover_size)));
                out_fifo_wr_en <= 1;
            end else if (unhandled_size > 0) begin
                if (leftover_size + unhandled_size >= AXI_WIDTH) begin
                    leftover_size <= leftover_size + unhandled_size - AXI_WIDTH;
                    leftover <= unhandled[curr] >> (AXI_WIDTH - leftover_size);
                    out_fifo_in <= (unhandled[curr] << leftover_size) + (leftover & (AXI_WIDTH'(-1) >> (AXI_WIDTH - leftover_size)));
                    out_fifo_wr_en <= 1;
                end else begin
                    leftover_size <= leftover_size + unhandled_size;
                    leftover <= (unhandled[curr] << leftover_size) | (leftover & (AXI_WIDTH'(-1) >> (AXI_WIDTH - leftover_size)));
                    out_fifo_wr_en <= 0;
                end
            end else if (do_finish && in_fifo_empty && ~din_valid) begin
                if (leftover_size > 0) begin
                    out_fifo_wr_en <= 1;
                    out_fifo_in <= leftover;
                    do_finish <= 0;
                end
            end else begin
                out_fifo_wr_en <= 0;
            end
`endif
        end
    end

    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            din_ready <= 0;
        end else begin
            din_ready <= ~in_fifo_almfull && ~out_fifo_almfull;
        end
    end

    logic [AXI_ADDR_WIDTH-1:0] buf_curr;
    logic [AXI_ADDR_WIDTH-1:0] buf_end;
    logic buf_write_en, buf_write_success;
    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            buf_curr <= 0;
            buf_end <= 0;
        end else if (buf_update) begin
            buf_curr <= buf_addr;
            buf_end <= buf_addr + buf_size;
        end else if (buf_write_en) begin
            buf_curr <= buf_curr + AXI_WIDTH/8;
        end

        interrupt <= (buf_curr == buf_end);
    end

    logic axi_aw_transmitted, axi_w_transmitted, axi_transmitted;
    logic axi_aw_working, axi_w_working, axi_working;
    assign axi_aw_transmitted = axi_out.awready & axi_out.awvalid;
    assign axi_w_transmitted = axi_out.wready & axi_out.wvalid;
    assign axi_aw_working = axi_out.awvalid & ~axi_out.awready;
    assign axi_w_working = axi_out.wvalid & ~axi_out.wready;
    assign axi_working = axi_aw_working | axi_w_working;

    // Transaction control
    logic axi_aw_handled, axi_w_handled;
    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            axi_aw_handled <= 0;
            axi_w_handled <= 0;
        end else begin
            if (axi_aw_transmitted & axi_w_transmitted) begin
                axi_aw_handled <= 0;
            end else if (axi_aw_transmitted) begin
                axi_aw_handled <= 1;
            end else if (axi_aw_handled & axi_w_transmitted) begin
                axi_aw_handled <= 0;
            end

            if (axi_aw_transmitted & axi_w_transmitted) begin
                axi_w_handled <= 0;
            end else if (axi_w_transmitted) begin
                axi_w_handled <= 1;
            end else if (axi_w_handled & axi_aw_handled) begin
                axi_w_handled <= 0;
            end
        end
    end

    assign axi_transmitted = (axi_aw_transmitted | axi_aw_handled) & (axi_w_transmitted | axi_w_handled);
    assign buf_write_en = axi_transmitted;

    // Valid control
    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            axi_out.awvalid <= 0;
            axi_out.wvalid <= 0;
        end else begin
            if (axi_aw_working) begin
                axi_out.awvalid <= 1;
            end else if (axi_w_working) begin
                axi_out.awvalid <= 0;
            end else begin
                axi_out.awvalid <= ~out_fifo_empty;
            end

            if (axi_w_working) begin
                axi_out.wvalid <= 1;
            end else if (axi_aw_working) begin
                axi_out.wvalid <= 0;
            end else begin
                axi_out.wvalid <= ~out_fifo_empty;
            end
        end
    end

    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            axi_out.wdata <= 0;
        end else begin
            if (~axi_aw_working & ~axi_w_working & ~out_fifo_empty)
                axi_out.wdata <= out_fifo_out;
        end
    end
    assign out_fifo_rd_en = ~axi_aw_working & ~axi_w_working & ~out_fifo_empty;

    logic [15:0] tid;
    always_ff @(posedge clk) begin
        if (~sync_rst_n) begin
            tid <= 0;
        end else begin
            if (axi_transmitted) begin
                tid <= tid + 1;
            end
        end
    end

    // AW extras
    assign axi_out.awid = tid;
    assign axi_out.awaddr = buf_curr;
    assign axi_out.awlen = 0;
    assign axi_out.awsize = AXI_WIDTH / 8;

    assign axi_out.wid = tid;
    assign axi_out.wstrb = -1;
    assign axi_out.wlast = 1;

    // Read and write response are always ready
    assign axi_out.bready = 1;
    assign axi_out.rready = 1;
endmodule
